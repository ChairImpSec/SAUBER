library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package emulate_bitstream is
--X0Y1, W_IO_custom
constant Tile_X0Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y1, linear_LMDPL
constant Tile_X1Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000000000000000000000";
--X2Y1, linear_LMDPL
constant Tile_X2Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010110101010101010100100010001000100000000000000000000100010001000100000000000000000";
--X3Y1, nonlinear_LMDPL
constant Tile_X3Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X4Y1, linear_LMDPL
constant Tile_X4Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X5Y1, linear_LMDPL
constant Tile_X5Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000000000001101110111011101000000000000000001000100010001000000000000000000";
--X6Y1, nonlinear_LMDPL
constant Tile_X6Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X7Y1, linear_LMDPL
constant Tile_X7Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110011011101110111010000000000000000";
--X8Y1, linear_LMDPL
constant Tile_X8Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100";
--X9Y1, nonlinear_LMDPL
constant Tile_X9Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X10Y1, linear_LMDPL
constant Tile_X10Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010001000100010000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X11Y1, linear_LMDPL
constant Tile_X11Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000100010001000100000000000000000000101010101010101";
--X12Y1, nonlinear_LMDPL
constant Tile_X12Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000001000100010001";
--X13Y1, linear_LMDPL
constant Tile_X13Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X14Y1, linear_LMDPL
constant Tile_X14Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X15Y1, nonlinear_LMDPL
constant Tile_X15Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000010001000100010000000000000000";
--X16Y1, linear_LMDPL
constant Tile_X16Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X17Y1, linear_LMDPL
constant Tile_X17Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X18Y1, nonlinear_LMDPL
constant Tile_X18Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001000100010001000";
--X19Y1, linear_LMDPL
constant Tile_X19Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X20Y1, linear_LMDPL
constant Tile_X20Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X21Y1, nonlinear_LMDPL
constant Tile_X21Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X22Y1, linear_LMDPL
constant Tile_X22Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X23Y1, linear_LMDPL
constant Tile_X23Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X24Y1, nonlinear_LMDPL
constant Tile_X24Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X25Y1, linear_LMDPL
constant Tile_X25Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X26Y1, linear_LMDPL
constant Tile_X26Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X27Y1, nonlinear_LMDPL
constant Tile_X27Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X28Y1, linear_LMDPL
constant Tile_X28Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001111111111111111";
--X29Y1, linear_LMDPL
constant Tile_X29Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000101010100000000000000000110011001100110001010101010101010000000000000000";
--X30Y1, nonlinear_LMDPL
constant Tile_X30Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y1, linear_LMDPL
constant Tile_X31Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001010101010101010";
--X32Y1, linear_LMDPL
constant Tile_X32Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000010101010000000000000000000000000101110111011101100000000000000001110111011101110";
--X33Y1, nonlinear_LMDPL
constant Tile_X33Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000000000000000000000";
--X34Y1, linear_LMDPL
constant Tile_X34Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X35Y1, linear_LMDPL
constant Tile_X35Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X36Y1, nonlinear_LMDPL
constant Tile_X36Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000010001000100010";
--X37Y1, linear_LMDPL
constant Tile_X37Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X38Y1, linear_LMDPL
constant Tile_X38Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X39Y1, nonlinear_LMDPL
constant Tile_X39Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X40Y1, linear_LMDPL
constant Tile_X40Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X41Y1, linear_LMDPL
constant Tile_X41Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010001000100010000000000000000000000000000000000011001100110011000000000000000000000000000000000";
--X42Y1, nonlinear_LMDPL
constant Tile_X42Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000001010101010101010000000000000000000000000010001000100010000000000101010100000000000000000100010001000100011111111111111110000000000000000";
--X43Y1, linear_LMDPL
constant Tile_X43Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000001100110011001101010101010101010000000000000000";
--X44Y1, linear_LMDPL
constant Tile_X44Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X45Y1, nonlinear_LMDPL
constant Tile_X45Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X46Y1, linear_LMDPL
constant Tile_X46Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X47Y1, linear_LMDPL
constant Tile_X47Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X48Y1, nonlinear_LMDPL
constant Tile_X48Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000001100110011001100000000000000001001100110011001";
--X49Y1, linear_LMDPL
constant Tile_X49Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X50Y1, linear_LMDPL
constant Tile_X50Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010101010101010100000000000000000101010101010101000000000000000000100010001000100000000000000000";
--X51Y1, nonlinear_LMDPL
constant Tile_X51Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000000000000000000000000000000000000";
--X52Y1, linear_LMDPL
constant Tile_X52Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X53Y1, linear_LMDPL
constant Tile_X53Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X54Y1, nonlinear_LMDPL
constant Tile_X54Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X55Y1, linear_LMDPL
constant Tile_X55Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X56Y1, linear_LMDPL
constant Tile_X56Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001100110011001100";
--X57Y1, nonlinear_LMDPL
constant Tile_X57Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X58Y1, linear_LMDPL
constant Tile_X58Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X59Y1, linear_LMDPL
constant Tile_X59Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X60Y1, nonlinear_LMDPL
constant Tile_X60Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y1, linear_LMDPL
constant Tile_X61Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X62Y1, linear_LMDPL
constant Tile_X62Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000101110111011101100110011001100110000000000000000";
--X63Y1, nonlinear_LMDPL
constant Tile_X63Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X64Y1, linear_LMDPL
constant Tile_X64Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X65Y1, linear_LMDPL
constant Tile_X65Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001111111111111111";
--X66Y1, nonlinear_LMDPL
constant Tile_X66Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X67Y1, linear_LMDPL
constant Tile_X67Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X68Y1, linear_LMDPL
constant Tile_X68Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X69Y1, nonlinear_LMDPL
constant Tile_X69Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X70Y1, linear_LMDPL
constant Tile_X70Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000001000100010001";
--X71Y1, linear_LMDPL
constant Tile_X71Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X72Y1, nonlinear_LMDPL
constant Tile_X72Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001101110111011101";
--X73Y1, linear_LMDPL
constant Tile_X73Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X74Y1, linear_LMDPL
constant Tile_X74Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X75Y1, nonlinear_LMDPL
constant Tile_X75Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X76Y1, linear_LMDPL
constant Tile_X76Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X77Y1, linear_LMDPL
constant Tile_X77Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X78Y1, ctrl_to_sec
constant Tile_X78Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y1, combined_WDDL
constant Tile_X79Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y1, combined_WDDL
constant Tile_X80Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y1, ctrl_IO
constant Tile_X81Y1_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y2, W_IO_custom
constant Tile_X0Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000";
--X1Y2, linear_LMDPL
constant Tile_X1Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000000001000100010001";
--X2Y2, linear_LMDPL
constant Tile_X2Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100100010001000100010000000000000000";
--X3Y2, nonlinear_LMDPL
constant Tile_X3Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000001010101010101010";
--X4Y2, linear_LMDPL
constant Tile_X4Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X5Y2, linear_LMDPL
constant Tile_X5Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000111011101110111";
--X6Y2, nonlinear_LMDPL
constant Tile_X6Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000001011101110111011";
--X7Y2, linear_LMDPL
constant Tile_X7Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000000000000000000011111111010101010101010100000000101010100011001100110011000000000000000010011001100110010000000000000000";
--X8Y2, linear_LMDPL
constant Tile_X8Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110010001000100010000000000000000000";
--X9Y2, nonlinear_LMDPL
constant Tile_X9Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000001000100010001";
--X10Y2, linear_LMDPL
constant Tile_X10Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111011101110";
--X11Y2, linear_LMDPL
constant Tile_X11Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X12Y2, nonlinear_LMDPL
constant Tile_X12Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101101010100000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X13Y2, linear_LMDPL
constant Tile_X13Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000011001100110011";
--X14Y2, linear_LMDPL
constant Tile_X14Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000011101110111011100000000000000001010101010101010";
--X15Y2, nonlinear_LMDPL
constant Tile_X15Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X16Y2, linear_LMDPL
constant Tile_X16Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X17Y2, linear_LMDPL
constant Tile_X17Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000010101010101010100101010100000000000000000000000000000000000000000000000000000000000100010001000100000000010101011110111011101110000000000000000000000000000000001100110011001100";
--X18Y2, nonlinear_LMDPL
constant Tile_X18Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X19Y2, linear_LMDPL
constant Tile_X19Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X20Y2, linear_LMDPL
constant Tile_X20Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X21Y2, nonlinear_LMDPL
constant Tile_X21Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X22Y2, linear_LMDPL
constant Tile_X22Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001011101110111011";
--X23Y2, linear_LMDPL
constant Tile_X23Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010001000100010000000000101010100000000000000000101110111011101100000000000000000000000000000000";
--X24Y2, nonlinear_LMDPL
constant Tile_X24Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X25Y2, linear_LMDPL
constant Tile_X25Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000101010100000000010101010000000000000000010101010000000000000000000000000000000000000000011111111000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X26Y2, linear_LMDPL
constant Tile_X26Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001100110011001100000000000000000";
--X27Y2, nonlinear_LMDPL
constant Tile_X27Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000010101010111111110000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000010001000100010";
--X28Y2, linear_LMDPL
constant Tile_X28Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001111111111111111";
--X29Y2, linear_LMDPL
constant Tile_X29Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X30Y2, nonlinear_LMDPL
constant Tile_X30Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000101010100000000000000000100010001000100000100010001000100000000000000000";
--X31Y2, linear_LMDPL
constant Tile_X31Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001100110011001100";
--X32Y2, linear_LMDPL
constant Tile_X32Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000011101110111011100000000000000000";
--X33Y2, nonlinear_LMDPL
constant Tile_X33Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000011111111000000000000000000000000101010100000000000000000001100110011001100000000000000000100010001000100";
--X34Y2, linear_LMDPL
constant Tile_X34Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000010101010101010100000000000000001100110011001100000000000000000010111011101110110000000000000000";
--X35Y2, linear_LMDPL
constant Tile_X35Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010010001000100010011111111000000000000000000000000001100110011001101000100010001000000000000000000";
--X36Y2, nonlinear_LMDPL
constant Tile_X36Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000001010101010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X37Y2, linear_LMDPL
constant Tile_X37Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001110111011101110110000000000000000";
--X38Y2, linear_LMDPL
constant Tile_X38Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X39Y2, nonlinear_LMDPL
constant Tile_X39Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000000100010001000100";
--X40Y2, linear_LMDPL
constant Tile_X40Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X41Y2, linear_LMDPL
constant Tile_X41Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010101010101000000000000000000100010001000100";
--X42Y2, nonlinear_LMDPL
constant Tile_X42Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000001010101000000000000000001010101010101010000000000000000000000000010101010101010100000000101010100100010001000100000000000000000000010001000100010000000000000000";
--X43Y2, linear_LMDPL
constant Tile_X43Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X44Y2, linear_LMDPL
constant Tile_X44Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111010101010000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X45Y2, nonlinear_LMDPL
constant Tile_X45Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101011101110111011000000000000000000000000000000001010101010101010";
--X46Y2, linear_LMDPL
constant Tile_X46Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X47Y2, linear_LMDPL
constant Tile_X47Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X48Y2, nonlinear_LMDPL
constant Tile_X48Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111111010101000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000011001100110011";
--X49Y2, linear_LMDPL
constant Tile_X49Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100001110111011101110000000000000000";
--X50Y2, linear_LMDPL
constant Tile_X50Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000100010001000100010101010101010100000000000000000";
--X51Y2, nonlinear_LMDPL
constant Tile_X51Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110101010100000000000000001010101000000000000000001111111111111111000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X52Y2, linear_LMDPL
constant Tile_X52Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000010101010000000000000000010101010101010101111111100000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X53Y2, linear_LMDPL
constant Tile_X53Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111010101010000000000000000010101010101010100000000101010100101010101010101000000000000000001100110011001100000000000000000";
--X54Y2, nonlinear_LMDPL
constant Tile_X54Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X55Y2, linear_LMDPL
constant Tile_X55Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X56Y2, linear_LMDPL
constant Tile_X56Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001000100010001000";
--X57Y2, nonlinear_LMDPL
constant Tile_X57Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001011101110111011";
--X58Y2, linear_LMDPL
constant Tile_X58Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X59Y2, linear_LMDPL
constant Tile_X59Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000001010101000000000010101010101010100000000000000000010001000100010000000000000000001110111011101110000000000000000";
--X60Y2, nonlinear_LMDPL
constant Tile_X60Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001011101110111011";
--X61Y2, linear_LMDPL
constant Tile_X61Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X62Y2, linear_LMDPL
constant Tile_X62Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000111111110000000010101010010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X63Y2, nonlinear_LMDPL
constant Tile_X63Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000100010001000100000000000000000001101110111011101";
--X64Y2, linear_LMDPL
constant Tile_X64Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001101110111011101000000000000000000100010001000100000000000000000";
--X65Y2, linear_LMDPL
constant Tile_X65Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X66Y2, nonlinear_LMDPL
constant Tile_X66Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101011010101000000000010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X67Y2, linear_LMDPL
constant Tile_X67Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X68Y2, linear_LMDPL
constant Tile_X68Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X69Y2, nonlinear_LMDPL
constant Tile_X69Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X70Y2, linear_LMDPL
constant Tile_X70Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X71Y2, linear_LMDPL
constant Tile_X71Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X72Y2, nonlinear_LMDPL
constant Tile_X72Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000010001000100010000000000000000";
--X73Y2, linear_LMDPL
constant Tile_X73Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X74Y2, linear_LMDPL
constant Tile_X74Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X75Y2, nonlinear_LMDPL
constant Tile_X75Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000001101110111011101";
--X76Y2, linear_LMDPL
constant Tile_X76Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X77Y2, linear_LMDPL
constant Tile_X77Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X78Y2, ctrl_to_sec
constant Tile_X78Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y2, combined_WDDL
constant Tile_X79Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y2, combined_WDDL
constant Tile_X80Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000";
--X81Y2, ctrl_IO
constant Tile_X81Y2_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000";
--X0Y3, W_IO_custom
constant Tile_X0Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y3, linear_LMDPL
constant Tile_X1Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000100110011001100101000100010001000000000000000000";
--X2Y3, linear_LMDPL
constant Tile_X2Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101111101110111011100000000000000000";
--X3Y3, nonlinear_LMDPL
constant Tile_X3Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X4Y3, linear_LMDPL
constant Tile_X4Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X5Y3, linear_LMDPL
constant Tile_X5Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100010111011101110110000000000000000";
--X6Y3, nonlinear_LMDPL
constant Tile_X6Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X7Y3, linear_LMDPL
constant Tile_X7Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111110101010010101010101010100000000000000000100010001000100000000000000000010011001100110010000000000000000";
--X8Y3, linear_LMDPL
constant Tile_X8Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001001100110011001";
--X9Y3, nonlinear_LMDPL
constant Tile_X9Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X10Y3, linear_LMDPL
constant Tile_X10Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000111101110111011100000000000000000";
--X11Y3, linear_LMDPL
constant Tile_X11Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000001010101000000000000000000000000101010100000000000000000001000100010001000000000000000000111011101110111";
--X12Y3, nonlinear_LMDPL
constant Tile_X12Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000011001100110011";
--X13Y3, linear_LMDPL
constant Tile_X13Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000000110011001100110";
--X14Y3, linear_LMDPL
constant Tile_X14Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001011101110111011";
--X15Y3, nonlinear_LMDPL
constant Tile_X15Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010011001100110010000000000000000";
--X16Y3, linear_LMDPL
constant Tile_X16Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X17Y3, linear_LMDPL
constant Tile_X17Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001111111100000000000000000000000000000000000000001010101010101010010101011010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X18Y3, nonlinear_LMDPL
constant Tile_X18Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010101111111100000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X19Y3, linear_LMDPL
constant Tile_X19Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000110011001100110";
--X20Y3, linear_LMDPL
constant Tile_X20Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000011111111000000000000000000000000000000000101010100000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X21Y3, nonlinear_LMDPL
constant Tile_X21Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000001010101000000000101010100000000000000000010101010101010100000000000000000101010101010101000000000000000001000100010001000000000000000000";
--X22Y3, linear_LMDPL
constant Tile_X22Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111111111111000000000101010110101010000000001010101000000000000000000000000011111111010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X23Y3, linear_LMDPL
constant Tile_X23Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000010101010010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X24Y3, nonlinear_LMDPL
constant Tile_X24Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X25Y3, linear_LMDPL
constant Tile_X25Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X26Y3, linear_LMDPL
constant Tile_X26Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X27Y3, nonlinear_LMDPL
constant Tile_X27Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X28Y3, linear_LMDPL
constant Tile_X28Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000100010001000110101010000000000101010101010101000000000000000000000000000000001000100010001000";
--X29Y3, linear_LMDPL
constant Tile_X29Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001011101110111011";
--X30Y3, nonlinear_LMDPL
constant Tile_X30Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101011010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000101110111011101100000000000000001101110111011101";
--X31Y3, linear_LMDPL
constant Tile_X31Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101000000000101010100101010100000000000000001010101000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X32Y3, linear_LMDPL
constant Tile_X32Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000001010101101010101010101010101010000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000110011001100110000000000000000";
--X33Y3, nonlinear_LMDPL
constant Tile_X33Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000001010101010101010101010100000000101010101100110011001100000000000000000010101010101010100000000000000000";
--X34Y3, linear_LMDPL
constant Tile_X34Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000010001000100010010111011101110110000000000000000";
--X35Y3, linear_LMDPL
constant Tile_X35Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000011111111010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X36Y3, nonlinear_LMDPL
constant Tile_X36Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000011011101110111010000000000000000";
--X37Y3, linear_LMDPL
constant Tile_X37Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X38Y3, linear_LMDPL
constant Tile_X38Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000101010110101010000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001010101010101010";
--X39Y3, nonlinear_LMDPL
constant Tile_X39Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000011111111000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X40Y3, linear_LMDPL
constant Tile_X40Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000011001100110011000000000000000001010101010101010000000000000000";
--X41Y3, linear_LMDPL
constant Tile_X41Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000010101010000000010101010010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X42Y3, nonlinear_LMDPL
constant Tile_X42Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000111111110101010110101010000000000000000000000000010001000100010000000000101010100000000000000000100110011001100101010101010101010000000000000000";
--X43Y3, linear_LMDPL
constant Tile_X43Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010101010100000000000000001101110111011101000000000000000000100010001000100000000000000000";
--X44Y3, linear_LMDPL
constant Tile_X44Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000001010101111111110000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X45Y3, nonlinear_LMDPL
constant Tile_X45Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000111111110101010100000000000000000101010100000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X46Y3, linear_LMDPL
constant Tile_X46Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000001010101000000001010101011111111000000000000000000000000000000000000000000000000010101010000000001010101010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X47Y3, linear_LMDPL
constant Tile_X47Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X48Y3, nonlinear_LMDPL
constant Tile_X48Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111010101010101010100000000101010101011101110111011000000000000000011001100110011000000000000000000";
--X49Y3, linear_LMDPL
constant Tile_X49Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X50Y3, linear_LMDPL
constant Tile_X50Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101111111100000000000100010001000100000000000000000011001100110011000000000000000000000000000000001000100010001000";
--X51Y3, nonlinear_LMDPL
constant Tile_X51Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001111111100000000101010101010101000000000000000000000000000000000000000000000000010101010010101010101010100000000101010100011001100110011000000000000000001000100010001000000000000000000";
--X52Y3, linear_LMDPL
constant Tile_X52Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010101010100000000001010101101010100000000001010101000000000000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X53Y3, linear_LMDPL
constant Tile_X53Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X54Y3, nonlinear_LMDPL
constant Tile_X54Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000111111110000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001010101010101010";
--X55Y3, linear_LMDPL
constant Tile_X55Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X56Y3, linear_LMDPL
constant Tile_X56Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101111111110000000000000000101010100000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X57Y3, nonlinear_LMDPL
constant Tile_X57Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000101010100000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X58Y3, linear_LMDPL
constant Tile_X58Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000100010001000100";
--X59Y3, linear_LMDPL
constant Tile_X59Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101011111111100000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X60Y3, nonlinear_LMDPL
constant Tile_X60Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X61Y3, linear_LMDPL
constant Tile_X61Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010101111111100000000010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X62Y3, linear_LMDPL
constant Tile_X62Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000010101010000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X63Y3, nonlinear_LMDPL
constant Tile_X63Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101001010101101010100000000011111111000000001010101000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X64Y3, linear_LMDPL
constant Tile_X64Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X65Y3, linear_LMDPL
constant Tile_X65Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001110111011101110";
--X66Y3, nonlinear_LMDPL
constant Tile_X66Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X67Y3, linear_LMDPL
constant Tile_X67Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011";
--X68Y3, linear_LMDPL
constant Tile_X68Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X69Y3, nonlinear_LMDPL
constant Tile_X69Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X70Y3, linear_LMDPL
constant Tile_X70Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000010001000100010";
--X71Y3, linear_LMDPL
constant Tile_X71Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X72Y3, nonlinear_LMDPL
constant Tile_X72Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000001000100010001000000000000000000";
--X73Y3, linear_LMDPL
constant Tile_X73Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000011001100110011";
--X74Y3, linear_LMDPL
constant Tile_X74Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100101010100000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000001000100010001";
--X75Y3, nonlinear_LMDPL
constant Tile_X75Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X76Y3, linear_LMDPL
constant Tile_X76Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001101110111011101";
--X77Y3, linear_LMDPL
constant Tile_X77Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000011001100110011";
--X78Y3, ctrl_to_sec
constant Tile_X78Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y3, combined_WDDL
constant Tile_X79Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y3, combined_WDDL
constant Tile_X80Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y3, ctrl_IO
constant Tile_X81Y3_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y4, W_IO_custom
constant Tile_X0Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000";
--X1Y4, linear_LMDPL
constant Tile_X1Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X2Y4, linear_LMDPL
constant Tile_X2Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010010101010000000000000000000000000011001100110011000010001000100010000000000000000";
--X3Y4, nonlinear_LMDPL
constant Tile_X3Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000110011001100110";
--X4Y4, linear_LMDPL
constant Tile_X4Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X5Y4, linear_LMDPL
constant Tile_X5Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000101010100000000010101010000000001010101000000000000000000000000011111111000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X6Y4, nonlinear_LMDPL
constant Tile_X6Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001100110011001100";
--X7Y4, linear_LMDPL
constant Tile_X7Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010111111110000000000000000101010100000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X8Y4, linear_LMDPL
constant Tile_X8Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000100010001000100000000000000000110011001100110";
--X9Y4, nonlinear_LMDPL
constant Tile_X9Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000110011001100110";
--X10Y4, linear_LMDPL
constant Tile_X10Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000010001000100010";
--X11Y4, linear_LMDPL
constant Tile_X11Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000001111111100000000000000001010101011111111000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X12Y4, nonlinear_LMDPL
constant Tile_X12Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X13Y4, linear_LMDPL
constant Tile_X13Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000100010001000100000000000000000001011101110111011";
--X14Y4, linear_LMDPL
constant Tile_X14Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X15Y4, nonlinear_LMDPL
constant Tile_X15Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X16Y4, linear_LMDPL
constant Tile_X16Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101011010101000000000000000000000000000000000000000001010101011111111000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X17Y4, linear_LMDPL
constant Tile_X17Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010101010101011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000101110111011101101000100010001000000000000000000";
--X18Y4, nonlinear_LMDPL
constant Tile_X18Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111100000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X19Y4, linear_LMDPL
constant Tile_X19Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010111111110000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X20Y4, linear_LMDPL
constant Tile_X20Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X21Y4, nonlinear_LMDPL
constant Tile_X21Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101111111101010101010001000100010000000000010101010000000000000000001000100010001000000000000000000000000000000000";
--X22Y4, linear_LMDPL
constant Tile_X22Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000101010101010101001010101010101010000000000000000";
--X23Y4, linear_LMDPL
constant Tile_X23Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X24Y4, nonlinear_LMDPL
constant Tile_X24Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000011111111010101010000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X25Y4, linear_LMDPL
constant Tile_X25Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001110111011101110000000000000000";
--X26Y4, linear_LMDPL
constant Tile_X26Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000001010101001010101000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001101110111011101000000000000000000100010001000100000000000000000";
--X27Y4, nonlinear_LMDPL
constant Tile_X27Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000001000100010001";
--X28Y4, linear_LMDPL
constant Tile_X28Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100101010100000000101010100000000010101010111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X29Y4, linear_LMDPL
constant Tile_X29Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X30Y4, nonlinear_LMDPL
constant Tile_X30Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000001000100010001";
--X31Y4, linear_LMDPL
constant Tile_X31Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010101010101010101000000000101010101010101010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X32Y4, linear_LMDPL
constant Tile_X32Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110011111111111111110000000000000000";
--X33Y4, nonlinear_LMDPL
constant Tile_X33Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000001010101000000000000000000000000010101010010001000100010000000000101010100000000000000000101110111011101101000100010001000000000000000000";
--X34Y4, linear_LMDPL
constant Tile_X34Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X35Y4, linear_LMDPL
constant Tile_X35Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X36Y4, nonlinear_LMDPL
constant Tile_X36Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000000100010001000100";
--X37Y4, linear_LMDPL
constant Tile_X37Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001011101110111011";
--X38Y4, linear_LMDPL
constant Tile_X38Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000000000000000000";
--X39Y4, nonlinear_LMDPL
constant Tile_X39Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111110101010010101010101010100000000101010101001100110011001000000000000000001000100010001000000000000000000";
--X40Y4, linear_LMDPL
constant Tile_X40Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000110111011101110101000100010001000000000000000000";
--X41Y4, linear_LMDPL
constant Tile_X41Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000100010001000100";
--X42Y4, nonlinear_LMDPL
constant Tile_X42Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000001010101010101010000000001111111100000000010101010101010100000000101010101001100110011001000000000000000001010101010101010000000000000000";
--X43Y4, linear_LMDPL
constant Tile_X43Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X44Y4, linear_LMDPL
constant Tile_X44Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010110101010000000000000000000000000101010100000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001101110111011101";
--X45Y4, nonlinear_LMDPL
constant Tile_X45Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X46Y4, linear_LMDPL
constant Tile_X46Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010110101010010101010000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X47Y4, linear_LMDPL
constant Tile_X47Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X48Y4, nonlinear_LMDPL
constant Tile_X48Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000101110111011101100010001000100010000000000000000";
--X49Y4, linear_LMDPL
constant Tile_X49Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X50Y4, linear_LMDPL
constant Tile_X50Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010101010101000000000010001000100010000000000101010100000000000000000111011101110111010111011101110110000000000000000";
--X51Y4, nonlinear_LMDPL
constant Tile_X51Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100101010100000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000001100110011001110011001100110010000000000000000";
--X52Y4, linear_LMDPL
constant Tile_X52Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X53Y4, linear_LMDPL
constant Tile_X53Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000010101010000000001010101000000000010101010101010100000000101010101100110011001100000000000000000001000100010001000000000000000000";
--X54Y4, nonlinear_LMDPL
constant Tile_X54Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000001010101001010101101010100000000000000000000000000000000000000000101010100000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X55Y4, linear_LMDPL
constant Tile_X55Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000010101010000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X56Y4, linear_LMDPL
constant Tile_X56Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000101010111111111010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000000011001100110011";
--X57Y4, nonlinear_LMDPL
constant Tile_X57Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000100010001000100";
--X58Y4, linear_LMDPL
constant Tile_X58Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X59Y4, linear_LMDPL
constant Tile_X59Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101011111111010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X60Y4, nonlinear_LMDPL
constant Tile_X60Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y4, linear_LMDPL
constant Tile_X61Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000011111111101010100101010100000000010001000100010000000000000000000000000000000000100010001000100010111011101110110000000000000000";
--X62Y4, linear_LMDPL
constant Tile_X62Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000010101010010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X63Y4, nonlinear_LMDPL
constant Tile_X63Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001011101110111011";
--X64Y4, linear_LMDPL
constant Tile_X64Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000110011001100110000000000000000010101010101010100000000000000000";
--X65Y4, linear_LMDPL
constant Tile_X65Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000101010100000000101010100000000000000000111111110000000000000000101010100000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001101110111011101";
--X66Y4, nonlinear_LMDPL
constant Tile_X66Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000100010001000100";
--X67Y4, linear_LMDPL
constant Tile_X67Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000110011001100110";
--X68Y4, linear_LMDPL
constant Tile_X68Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X69Y4, nonlinear_LMDPL
constant Tile_X69Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X70Y4, linear_LMDPL
constant Tile_X70Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000001111111100000000010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X71Y4, linear_LMDPL
constant Tile_X71Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X72Y4, nonlinear_LMDPL
constant Tile_X72Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X73Y4, linear_LMDPL
constant Tile_X73Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000101010101010101";
--X74Y4, linear_LMDPL
constant Tile_X74Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X75Y4, nonlinear_LMDPL
constant Tile_X75Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000010001000100010";
--X76Y4, linear_LMDPL
constant Tile_X76Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X77Y4, linear_LMDPL
constant Tile_X77Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X78Y4, ctrl_to_sec
constant Tile_X78Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y4, combined_WDDL
constant Tile_X79Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y4, combined_WDDL
constant Tile_X80Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y4, ctrl_IO
constant Tile_X81Y4_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y5, W_IO_custom
constant Tile_X0Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000";
--X1Y5, linear_LMDPL
constant Tile_X1Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X2Y5, linear_LMDPL
constant Tile_X2Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000001000100010001";
--X3Y5, nonlinear_LMDPL
constant Tile_X3Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X4Y5, linear_LMDPL
constant Tile_X4Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X5Y5, linear_LMDPL
constant Tile_X5Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010110101010000100010001000100000000000000000011001100110011000000000000000000000000000000001001100110011001";
--X6Y5, nonlinear_LMDPL
constant Tile_X6Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X7Y5, linear_LMDPL
constant Tile_X7Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X8Y5, linear_LMDPL
constant Tile_X8Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000001000100010001";
--X9Y5, nonlinear_LMDPL
constant Tile_X9Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X10Y5, linear_LMDPL
constant Tile_X10Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X11Y5, linear_LMDPL
constant Tile_X11Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101001100110011001000000000000000011011101110111010000000000000000";
--X12Y5, nonlinear_LMDPL
constant Tile_X12Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000010001000100010000000000000000";
--X13Y5, linear_LMDPL
constant Tile_X13Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X14Y5, linear_LMDPL
constant Tile_X14Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000010101010101010101010101010101010000100010001000100000000000000000101010101010101000000000000000000000000000000001110111011101110";
--X15Y5, nonlinear_LMDPL
constant Tile_X15Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X16Y5, linear_LMDPL
constant Tile_X16Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100101010100000000000000001010101000000000000000000000000000000000000000001010101010101010010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X17Y5, linear_LMDPL
constant Tile_X17Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X18Y5, nonlinear_LMDPL
constant Tile_X18Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y5, linear_LMDPL
constant Tile_X19Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X20Y5, linear_LMDPL
constant Tile_X20Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X21Y5, nonlinear_LMDPL
constant Tile_X21Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X22Y5, linear_LMDPL
constant Tile_X22Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000101010100000000001010101000000001010101000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X23Y5, linear_LMDPL
constant Tile_X23Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000010101010000000010101010010101010101010100000000000000000111011101110111000000000000000000110011001100110000000000000000";
--X24Y5, nonlinear_LMDPL
constant Tile_X24Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X25Y5, linear_LMDPL
constant Tile_X25Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000001010101000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X26Y5, linear_LMDPL
constant Tile_X26Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000001111111100000000010101010101010100000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X27Y5, nonlinear_LMDPL
constant Tile_X27Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111010101010000000000000000101010100000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X28Y5, linear_LMDPL
constant Tile_X28Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101001010101000000000000000000000000111111110000000010101010000000000000000000000000010001000100010000000000000000000000000000000000111011101110111001010101010101010000000000000000";
--X29Y5, linear_LMDPL
constant Tile_X29Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010100100010001000100000000000000000000100010001000100000000000000000";
--X30Y5, nonlinear_LMDPL
constant Tile_X30Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X31Y5, linear_LMDPL
constant Tile_X31Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000010101010101010110101010000000000000000000000000101010101010101000000000010101010101010100000000000000001010101000000000000000000000000011111111010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X32Y5, linear_LMDPL
constant Tile_X32Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X33Y5, nonlinear_LMDPL
constant Tile_X33Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000000011001100110011";
--X34Y5, linear_LMDPL
constant Tile_X34Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X35Y5, linear_LMDPL
constant Tile_X35Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111111111110000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000001000100010001000";
--X36Y5, nonlinear_LMDPL
constant Tile_X36Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y5, linear_LMDPL
constant Tile_X37Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010011011101110111010000000000000000";
--X38Y5, linear_LMDPL
constant Tile_X38Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X39Y5, nonlinear_LMDPL
constant Tile_X39Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000011111111010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X40Y5, linear_LMDPL
constant Tile_X40Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101011111111000000000000000010101010000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X41Y5, linear_LMDPL
constant Tile_X41Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X42Y5, nonlinear_LMDPL
constant Tile_X42Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010001000100010000000000101010100000000000000000000000000000000010011001100110010000000000000000";
--X43Y5, linear_LMDPL
constant Tile_X43Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X44Y5, linear_LMDPL
constant Tile_X44Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X45Y5, nonlinear_LMDPL
constant Tile_X45Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000100010001000100";
--X46Y5, linear_LMDPL
constant Tile_X46Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000001010101000000000101010100000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101010101010101010100000000000000000";
--X47Y5, linear_LMDPL
constant Tile_X47Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X48Y5, nonlinear_LMDPL
constant Tile_X48Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000001000100010001000";
--X49Y5, linear_LMDPL
constant Tile_X49Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000101010101111111110101010010101010101010100000000010101011100110011001100000000000000000001000100010001000000000000000000";
--X50Y5, linear_LMDPL
constant Tile_X50Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000001010101101010100000000000000000000000000000000000000000000000000101010100000000000000001010101000000000101010101010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X51Y5, nonlinear_LMDPL
constant Tile_X51Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X52Y5, linear_LMDPL
constant Tile_X52Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000000000000101010100000000000000000000000001010101000000000000000010101010111111110000000000000000101010100101010100000000101010100000000010101010000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001100110011001100";
--X53Y5, linear_LMDPL
constant Tile_X53Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010101011111111100000000010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X54Y5, nonlinear_LMDPL
constant Tile_X54Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010101010101010100110011001100110000000000000000";
--X55Y5, linear_LMDPL
constant Tile_X55Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X56Y5, linear_LMDPL
constant Tile_X56Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X57Y5, nonlinear_LMDPL
constant Tile_X57Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X58Y5, linear_LMDPL
constant Tile_X58Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001111111100000000010101010000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X59Y5, linear_LMDPL
constant Tile_X59Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101011010101000000000010001000100010000000000000000000000000000000000101110111011101110101010101010100000000000000000";
--X60Y5, nonlinear_LMDPL
constant Tile_X60Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000001000100010001000";
--X61Y5, linear_LMDPL
constant Tile_X61Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000101010100000000000000000000000001010101000000000101010100000000001010101000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X62Y5, linear_LMDPL
constant Tile_X62Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000001010101000000000111111110101010110101010010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X63Y5, nonlinear_LMDPL
constant Tile_X63Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000001010101101010100000000010101010000000001010101000000000010101011010101010101010010001000100010000000000000000000000000000000000001100110011001100100010001000100000000000000000";
--X64Y5, linear_LMDPL
constant Tile_X64Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000010101010101010100000000101010100000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X65Y5, linear_LMDPL
constant Tile_X65Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000010001000100010";
--X66Y5, nonlinear_LMDPL
constant Tile_X66Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000101010101010101010001000100010000000000000000000000000000000000001100110011001100100010001000100000000000000000";
--X67Y5, linear_LMDPL
constant Tile_X67Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X68Y5, linear_LMDPL
constant Tile_X68Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X69Y5, nonlinear_LMDPL
constant Tile_X69Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X70Y5, linear_LMDPL
constant Tile_X70Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000100010001000100000000000000000000010001000100010";
--X71Y5, linear_LMDPL
constant Tile_X71Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000101010101010101000010001000100010000000000000000";
--X72Y5, nonlinear_LMDPL
constant Tile_X72Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001101110111011101";
--X73Y5, linear_LMDPL
constant Tile_X73Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X74Y5, linear_LMDPL
constant Tile_X74Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000001010101001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X75Y5, nonlinear_LMDPL
constant Tile_X75Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X76Y5, linear_LMDPL
constant Tile_X76Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X77Y5, linear_LMDPL
constant Tile_X77Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000101100110011001100000000000000000";
--X78Y5, ctrl_to_sec
constant Tile_X78Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y5, combined_WDDL
constant Tile_X79Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y5, combined_WDDL
constant Tile_X80Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y5, ctrl_IO
constant Tile_X81Y5_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000";
--X0Y6, W_IO_custom
constant Tile_X0Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000111111110000000000000000000000000000000010100000000000000000000000000000000";
--X1Y6, linear_LMDPL
constant Tile_X1Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101100010001000100010000000000000000";
--X2Y6, linear_LMDPL
constant Tile_X2Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010100000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X3Y6, nonlinear_LMDPL
constant Tile_X3Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000010001000100010";
--X4Y6, linear_LMDPL
constant Tile_X4Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001000100010001000";
--X5Y6, linear_LMDPL
constant Tile_X5Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X6Y6, nonlinear_LMDPL
constant Tile_X6Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001001100110011001";
--X7Y6, linear_LMDPL
constant Tile_X7Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001111111111111111";
--X8Y6, linear_LMDPL
constant Tile_X8Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000100010001000100";
--X9Y6, nonlinear_LMDPL
constant Tile_X9Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000100110011001100100000000000000001010101010101010";
--X10Y6, linear_LMDPL
constant Tile_X10Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X11Y6, linear_LMDPL
constant Tile_X11Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001100110011001100";
--X12Y6, nonlinear_LMDPL
constant Tile_X12Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000001000100010001000000000000000010001000100010000000000000000000";
--X13Y6, linear_LMDPL
constant Tile_X13Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010011101110111011100000000000000000";
--X14Y6, linear_LMDPL
constant Tile_X14Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000010101010101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000111111111111111110101010101010100000000000000000";
--X15Y6, nonlinear_LMDPL
constant Tile_X15Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010001000100010000000000010101010000000000000000100110011001100110001000100010000000000000000000";
--X16Y6, linear_LMDPL
constant Tile_X16Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X17Y6, linear_LMDPL
constant Tile_X17Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000001000100010001000";
--X18Y6, nonlinear_LMDPL
constant Tile_X18Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101110111011101110011001100110010000000000000000";
--X19Y6, linear_LMDPL
constant Tile_X19Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000011001100110011";
--X20Y6, linear_LMDPL
constant Tile_X20Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X21Y6, nonlinear_LMDPL
constant Tile_X21Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000100010001000100000000101010101001100110011001000000000000000000000000000000001101110111011101";
--X22Y6, linear_LMDPL
constant Tile_X22Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000010101010000000000000000010101010101010100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X23Y6, linear_LMDPL
constant Tile_X23Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000001010101010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X24Y6, nonlinear_LMDPL
constant Tile_X24Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000011111111000000001010101010101010000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000011001100110011001000100010001000000000000000000";
--X25Y6, linear_LMDPL
constant Tile_X25Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000110011001100110000000000000000";
--X26Y6, linear_LMDPL
constant Tile_X26Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X27Y6, nonlinear_LMDPL
constant Tile_X27Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000010101010101010100101010101010101000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X28Y6, linear_LMDPL
constant Tile_X28Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010010101010000000000000000000000000100010001000100001100110011001100000000000000000";
--X29Y6, linear_LMDPL
constant Tile_X29Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000101010101010101011111111000000000000000000000000000000000000000011111111000000001111111100000000010001000100010000000000010101010000000000000000111111111111111101000100010001000000000000000000";
--X30Y6, nonlinear_LMDPL
constant Tile_X30Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000101010100000000000000000001100110011001100110011001100110000000000000000";
--X31Y6, linear_LMDPL
constant Tile_X31Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101011010101010101010000000000000000011111111000000001010101011111111010101010101010100000000000000001010101010101010111111110000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X32Y6, linear_LMDPL
constant Tile_X32Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000011111111101010101010101010101010000000000000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X33Y6, nonlinear_LMDPL
constant Tile_X33Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000001010101000000000010101010000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000000011001100110011";
--X34Y6, linear_LMDPL
constant Tile_X34Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000110111011101110100000000000000001100110011001100";
--X35Y6, linear_LMDPL
constant Tile_X35Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001011101110111011";
--X36Y6, nonlinear_LMDPL
constant Tile_X36Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y6, linear_LMDPL
constant Tile_X37Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X38Y6, linear_LMDPL
constant Tile_X38Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X39Y6, nonlinear_LMDPL
constant Tile_X39Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000101110111011101110001000100010000000000000000000";
--X40Y6, linear_LMDPL
constant Tile_X40Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X41Y6, linear_LMDPL
constant Tile_X41Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000010101010000100010001000100000000101010100011001100110011000000000000000000000000000000000010001000100010";
--X42Y6, nonlinear_LMDPL
constant Tile_X42Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111010101010101010100000000101010101100110011001100000000000000000010111011101110110000000000000000";
--X43Y6, linear_LMDPL
constant Tile_X43Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X44Y6, linear_LMDPL
constant Tile_X44Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X45Y6, nonlinear_LMDPL
constant Tile_X45Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000000000000000000010011001100110010000000000000000";
--X46Y6, linear_LMDPL
constant Tile_X46Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X47Y6, linear_LMDPL
constant Tile_X47Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X48Y6, nonlinear_LMDPL
constant Tile_X48Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000101010100001000100010001000000000000000001000100010001000000000000000000";
--X49Y6, linear_LMDPL
constant Tile_X49Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111010101011010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X50Y6, linear_LMDPL
constant Tile_X50Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010101010000000000000000000000001010101000000000000000001010101000000000000000000101010100000000000000001010101000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X51Y6, nonlinear_LMDPL
constant Tile_X51Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100101010101010101000000001010101000000000010101010000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X52Y6, linear_LMDPL
constant Tile_X52Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000101010110101010010101010000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X53Y6, linear_LMDPL
constant Tile_X53Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010101111111101010101010101010101010100000000101010101101110111011101000000000000000010001000100010000000000000000000";
--X54Y6, nonlinear_LMDPL
constant Tile_X54Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000001010101000000000101010100000000000000000000000001010101000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X55Y6, linear_LMDPL
constant Tile_X55Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010111111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X56Y6, linear_LMDPL
constant Tile_X56Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001100110011001100";
--X57Y6, nonlinear_LMDPL
constant Tile_X57Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000010101010000000000000000000000000000000011111111000000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000101010101010101";
--X58Y6, linear_LMDPL
constant Tile_X58Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101101010100000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X59Y6, linear_LMDPL
constant Tile_X59Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000010101010101010101010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X60Y6, nonlinear_LMDPL
constant Tile_X60Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000010101010000000001010101010101010101010100000000101010100100010001000100000000000000000000110011001100110000000000000000";
--X61Y6, linear_LMDPL
constant Tile_X61Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000010101010101010100000000010101010000000000000000010101010101010100101010100000000000100010001000100000000000000001011101110111011000000000000000000000000000000001100110011001100";
--X62Y6, linear_LMDPL
constant Tile_X62Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000100010001000100010111011101110110000000000000000";
--X63Y6, nonlinear_LMDPL
constant Tile_X63Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100000000010101010000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000001000100010001000000000000000000100010001000100";
--X64Y6, linear_LMDPL
constant Tile_X64Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X65Y6, linear_LMDPL
constant Tile_X65Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000101010100000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111111111111111100110011001100110000000000000000";
--X66Y6, nonlinear_LMDPL
constant Tile_X66Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101011011101110111011000000000000000010101010101010100000000000000000";
--X67Y6, linear_LMDPL
constant Tile_X67Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X68Y6, linear_LMDPL
constant Tile_X68Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X69Y6, nonlinear_LMDPL
constant Tile_X69Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X70Y6, linear_LMDPL
constant Tile_X70Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101";
--X71Y6, linear_LMDPL
constant Tile_X71Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X72Y6, nonlinear_LMDPL
constant Tile_X72Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X73Y6, linear_LMDPL
constant Tile_X73Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X74Y6, linear_LMDPL
constant Tile_X74Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X75Y6, nonlinear_LMDPL
constant Tile_X75Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X76Y6, linear_LMDPL
constant Tile_X76Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000100010001000100000000000000001101110111011101000000000000000000000000000000000101010101010101";
--X77Y6, linear_LMDPL
constant Tile_X77Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000101010101010101";
--X78Y6, ctrl_to_sec
constant Tile_X78Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y6, combined_WDDL
constant Tile_X79Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y6, combined_WDDL
constant Tile_X80Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y6, ctrl_IO
constant Tile_X81Y6_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000000";
--X0Y7, W_IO_custom
constant Tile_X0Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000001111111100000000010000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000";
--X1Y7, linear_LMDPL
constant Tile_X1Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X2Y7, linear_LMDPL
constant Tile_X2Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000100010001000100000000000000000010111011101110110000000000000000";
--X3Y7, nonlinear_LMDPL
constant Tile_X3Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001010101010101010";
--X4Y7, linear_LMDPL
constant Tile_X4Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X5Y7, linear_LMDPL
constant Tile_X5Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X6Y7, nonlinear_LMDPL
constant Tile_X6Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X7Y7, linear_LMDPL
constant Tile_X7Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000011111111000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X8Y7, linear_LMDPL
constant Tile_X8Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000100010001000110101010000000001100110011001100000000000000000000000000000000000011001100110011";
--X9Y7, nonlinear_LMDPL
constant Tile_X9Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000001010101000000000101010101010101011111111000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X10Y7, linear_LMDPL
constant Tile_X10Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000001010101000000001010101000000000101010100000000000000000000000000101010100000000000000000000000010101010010001000100010000000000000000000000000000000000111111111111111100100010001000100000000000000000";
--X11Y7, linear_LMDPL
constant Tile_X11Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000101010100011001100110011000000000000000001000100010001000000000000000000";
--X12Y7, nonlinear_LMDPL
constant Tile_X12Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X13Y7, linear_LMDPL
constant Tile_X13Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X14Y7, linear_LMDPL
constant Tile_X14Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000010101010101010100000000010101010000000001111111110101010101010100000000011111111010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X15Y7, nonlinear_LMDPL
constant Tile_X15Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000010101010101010100000000000000001001100110011001000000000000000011001100110011000000000000000000";
--X16Y7, linear_LMDPL
constant Tile_X16Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000011101110111011100000000000000001010101010101010";
--X17Y7, linear_LMDPL
constant Tile_X17Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000101010100000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X18Y7, nonlinear_LMDPL
constant Tile_X18Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001100110011001100010001000100010000000000000000";
--X19Y7, linear_LMDPL
constant Tile_X19Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X20Y7, linear_LMDPL
constant Tile_X20Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X21Y7, nonlinear_LMDPL
constant Tile_X21Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010001000100010000000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X22Y7, linear_LMDPL
constant Tile_X22Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000001010101000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001111111111111111";
--X23Y7, linear_LMDPL
constant Tile_X23Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X24Y7, nonlinear_LMDPL
constant Tile_X24Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000001000100010001010001000100010000000000000000000";
--X25Y7, linear_LMDPL
constant Tile_X25Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X26Y7, linear_LMDPL
constant Tile_X26Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100101010111111111000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X27Y7, nonlinear_LMDPL
constant Tile_X27Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000001010101010101010101010101010101010101010000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X28Y7, linear_LMDPL
constant Tile_X28Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000101010100000000111111111010101010101010000000001010101000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X29Y7, linear_LMDPL
constant Tile_X29Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010010101010000000001010101000000000000000010101010000000001010101011111111010001000100010000000000101010100000000000000000101010101010101011011101110111010000000000000000";
--X30Y7, nonlinear_LMDPL
constant Tile_X30Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101000000000000000000000000000000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000001100110011001111011101110111010000000000000000";
--X31Y7, linear_LMDPL
constant Tile_X31Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111101010101101010100000000000000000000000000000000000000000000000000000000001010101010101010000000000000000101010101010101011111111000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X32Y7, linear_LMDPL
constant Tile_X32Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111111111111000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001010101010101010";
--X33Y7, nonlinear_LMDPL
constant Tile_X33Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000010101010000000001010101000000000101010100000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000000010001000100010";
--X34Y7, linear_LMDPL
constant Tile_X34Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X35Y7, linear_LMDPL
constant Tile_X35Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X36Y7, nonlinear_LMDPL
constant Tile_X36Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100100010001000100000000000000000000000000000000000011001100110011";
--X37Y7, linear_LMDPL
constant Tile_X37Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X38Y7, linear_LMDPL
constant Tile_X38Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000010101011111111100000000010101010101010100000000010101010010001000100010000000000000000001000100010001000000000000000000";
--X39Y7, nonlinear_LMDPL
constant Tile_X39Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X40Y7, linear_LMDPL
constant Tile_X40Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100101010100000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000110111011101110110111011101110110000000000000000";
--X41Y7, linear_LMDPL
constant Tile_X41Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X42Y7, nonlinear_LMDPL
constant Tile_X42Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000100010001000100";
--X43Y7, linear_LMDPL
constant Tile_X43Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X44Y7, linear_LMDPL
constant Tile_X44Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X45Y7, nonlinear_LMDPL
constant Tile_X45Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000011011101110111010000000000000000";
--X46Y7, linear_LMDPL
constant Tile_X46Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011111111100000000000000000101010100000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010111111111000000001010101000000000101010100000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001101110111011101";
--X47Y7, linear_LMDPL
constant Tile_X47Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101010101010000000000000000011111111000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X48Y7, nonlinear_LMDPL
constant Tile_X48Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010110101010000000000000000000000000101010100000000000000000100010001000100000000000000000001001100110011001";
--X49Y7, linear_LMDPL
constant Tile_X49Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000111111111010101000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X50Y7, linear_LMDPL
constant Tile_X50Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000001010101000000000000000000000000001010101000000000101010100000000000000001010101000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X51Y7, nonlinear_LMDPL
constant Tile_X51Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101011111111100000000000000000000000001010101000000001010101001010101101010100000000001010101000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001000100010001000000000000000000001010101010101010000000000000000";
--X52Y7, linear_LMDPL
constant Tile_X52Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000010101011010101000000000111111110000000010101010000000001010101000000000000000000000000001010101010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X53Y7, linear_LMDPL
constant Tile_X53Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000000000001111111100000000010101010000000000000000000000000101010100000000000000000000000010101010000000001010101000000000000000000000000010101010010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X54Y7, nonlinear_LMDPL
constant Tile_X54Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X55Y7, linear_LMDPL
constant Tile_X55Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000111111110000000001010101000000000000000000000000101010100000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001111111111111111";
--X56Y7, linear_LMDPL
constant Tile_X56Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101111111110000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X57Y7, nonlinear_LMDPL
constant Tile_X57Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110";
--X58Y7, linear_LMDPL
constant Tile_X58Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000001010101101010100000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000110011001100110000000000000000001000100010001000";
--X59Y7, linear_LMDPL
constant Tile_X59Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000001010101000000000101010100000000101010101111111100000000010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X60Y7, nonlinear_LMDPL
constant Tile_X60Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000011111111000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X61Y7, linear_LMDPL
constant Tile_X61Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000101010111111111010101010000000010101010000000000000000000000000101010100000000001010101000100010001000100000000000000000101010101010101000000000000000000000000000000001011101110111011";
--X62Y7, linear_LMDPL
constant Tile_X62Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X63Y7, nonlinear_LMDPL
constant Tile_X63Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000001010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X64Y7, linear_LMDPL
constant Tile_X64Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000010101010000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X65Y7, linear_LMDPL
constant Tile_X65Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X66Y7, nonlinear_LMDPL
constant Tile_X66Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X67Y7, linear_LMDPL
constant Tile_X67Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X68Y7, linear_LMDPL
constant Tile_X68Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X69Y7, nonlinear_LMDPL
constant Tile_X69Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X70Y7, linear_LMDPL
constant Tile_X70Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010010101010000000001010101000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000101010101010101011101110111011100000000000000000";
--X71Y7, linear_LMDPL
constant Tile_X71Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X72Y7, nonlinear_LMDPL
constant Tile_X72Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X73Y7, linear_LMDPL
constant Tile_X73Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000011011101110111010000000000000000";
--X74Y7, linear_LMDPL
constant Tile_X74Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X75Y7, nonlinear_LMDPL
constant Tile_X75Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000101010100000000000000000010101010101010100000000111111111011101110111011000000000000000000010001000100010000000000000000";
--X76Y7, linear_LMDPL
constant Tile_X76Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000011001100110011";
--X77Y7, linear_LMDPL
constant Tile_X77Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000101010101000000000101010101010101000000000000000000000000000000000000000000000000";
--X78Y7, ctrl_to_sec
constant Tile_X78Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y7, combined_WDDL
constant Tile_X79Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y7, combined_WDDL
constant Tile_X80Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y7, ctrl_IO
constant Tile_X81Y7_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y8, W_IO_custom
constant Tile_X0Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000";
--X1Y8, linear_LMDPL
constant Tile_X1Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000001100110011001100000000000000000";
--X2Y8, linear_LMDPL
constant Tile_X2Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000001010101000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X3Y8, nonlinear_LMDPL
constant Tile_X3Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000001010101101010100000000001010101000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000011101110111011100000000000000001100110011001100";
--X4Y8, linear_LMDPL
constant Tile_X4Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X5Y8, linear_LMDPL
constant Tile_X5Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000011001100110011000000000000000001100110011001100";
--X6Y8, nonlinear_LMDPL
constant Tile_X6Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000010101010010001000100010000000000000000000000000000000000010001000100010";
--X7Y8, linear_LMDPL
constant Tile_X7Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X8Y8, linear_LMDPL
constant Tile_X8Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101010101010101010100000000101010100000000000000000000000000000000000010001000100010000000000000000";
--X9Y8, nonlinear_LMDPL
constant Tile_X9Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000001010101000000001010101000000000101010100000000000000000000000001010101000000000101010100000000001010101000000000000000000000000000000001010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000010001000100010";
--X10Y8, linear_LMDPL
constant Tile_X10Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010111111111000000001010101000000000111111110000000000000000000000001010101010101010000000000000000010101010010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X11Y8, linear_LMDPL
constant Tile_X11Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010101010101010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000110011001100110";
--X12Y8, nonlinear_LMDPL
constant Tile_X12Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X13Y8, linear_LMDPL
constant Tile_X13Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X14Y8, linear_LMDPL
constant Tile_X14Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000010101010101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100110011001100110101010101010100000000000000000";
--X15Y8, nonlinear_LMDPL
constant Tile_X15Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110010111011101110110000000000000000";
--X16Y8, linear_LMDPL
constant Tile_X16Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000001010101011111111000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X17Y8, linear_LMDPL
constant Tile_X17Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X18Y8, nonlinear_LMDPL
constant Tile_X18Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010111111111000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001001100110011001";
--X19Y8, linear_LMDPL
constant Tile_X19Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010110101010101010100000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000011101110111011100000000000000001000100010001000";
--X20Y8, linear_LMDPL
constant Tile_X20Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000100010001000100000000000000000001110111011101110000000000000000";
--X21Y8, nonlinear_LMDPL
constant Tile_X21Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000101010100000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000000000000011001100110011000000000000000000001000100010001";
--X22Y8, linear_LMDPL
constant Tile_X22Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000111111110000000001010101010101010101010100000000101010100000000000000000000000000000000000110011001100110000000000000000";
--X23Y8, linear_LMDPL
constant Tile_X23Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X24Y8, nonlinear_LMDPL
constant Tile_X24Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X25Y8, linear_LMDPL
constant Tile_X25Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000001100110011001100";
--X26Y8, linear_LMDPL
constant Tile_X26Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010101111111110101010010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X27Y8, nonlinear_LMDPL
constant Tile_X27Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101010101010101010100101010100000000000000000000000000000000000000000000000010101010010101010101010100000000000000001011101110111011000000000000000001010101010101010000000000000000";
--X28Y8, linear_LMDPL
constant Tile_X28Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101011111111000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X29Y8, linear_LMDPL
constant Tile_X29Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000001010101000000000000000000101010100000000101010100000000010101010101010101010101010101010010101010000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X30Y8, nonlinear_LMDPL
constant Tile_X30Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000101010101011101110111011000000000000000001000100010001000000000000000000";
--X31Y8, linear_LMDPL
constant Tile_X31Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001110111011101110";
--X32Y8, linear_LMDPL
constant Tile_X32Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000101010101010101010101010010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000111011101110111000000000000000001000100010001000000000000000000";
--X33Y8, nonlinear_LMDPL
constant Tile_X33Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000101010100000000010101010000000000000000000000001010101010101010000000000000000000000000000000000101010100000000000000000000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000001110111011101110";
--X34Y8, linear_LMDPL
constant Tile_X34Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X35Y8, linear_LMDPL
constant Tile_X35Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000011111111000000000101010100000000000000000000000010101010010101010101010100000000000000001111111111111111000000000000000000100010001000100000000000000000";
--X36Y8, nonlinear_LMDPL
constant Tile_X36Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y8, linear_LMDPL
constant Tile_X37Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000001010101101010101010101000000000101010100000000000000000000000000000000000000000101010100000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X38Y8, linear_LMDPL
constant Tile_X38Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111111010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000001010101000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001101110111011101";
--X39Y8, nonlinear_LMDPL
constant Tile_X39Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X40Y8, linear_LMDPL
constant Tile_X40Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000011001100110011";
--X41Y8, linear_LMDPL
constant Tile_X41Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000010101010010101010101010100000000101010100100010001000100000000000000000001010101010101010000000000000000";
--X42Y8, nonlinear_LMDPL
constant Tile_X42Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000011111111010101010101010100000000101010100000000000000000000000000000000010011001100110010000000000000000";
--X43Y8, linear_LMDPL
constant Tile_X43Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X44Y8, linear_LMDPL
constant Tile_X44Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000001000100010001000000000000000000101010101010101";
--X45Y8, nonlinear_LMDPL
constant Tile_X45Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011";
--X46Y8, linear_LMDPL
constant Tile_X46Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000001010101000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X47Y8, linear_LMDPL
constant Tile_X47Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000001010101010101010101010100000000010101010000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X48Y8, nonlinear_LMDPL
constant Tile_X48Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000001010101010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000010001000100010";
--X49Y8, linear_LMDPL
constant Tile_X49Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000111111110101010100000000010101010101010100000000000000000111011101110111000000000000000011001100110011000000000000000000";
--X50Y8, linear_LMDPL
constant Tile_X50Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010101010101000000000000000000000000000000001010101000000000010101010101010100000000101010100010001000100010000000000000000010001000100010000000000000000000";
--X51Y8, nonlinear_LMDPL
constant Tile_X51Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001111111100000000000000001010101000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X52Y8, linear_LMDPL
constant Tile_X52Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000001010101000000000101010100000000010101010101010100000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000010101010101010100000000000000000";
--X53Y8, linear_LMDPL
constant Tile_X53Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111111111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010101010101000000000000000000011001100110011";
--X54Y8, nonlinear_LMDPL
constant Tile_X54Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000101010101010101000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X55Y8, linear_LMDPL
constant Tile_X55Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X56Y8, linear_LMDPL
constant Tile_X56Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000001111111100000000101010100101010100000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000100010001000100001000100010001000000000000000000";
--X57Y8, nonlinear_LMDPL
constant Tile_X57Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010110101010010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000010001000100010";
--X58Y8, linear_LMDPL
constant Tile_X58Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X59Y8, linear_LMDPL
constant Tile_X59Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000010101010000000000000000010101010101010101010101000000000010101010101010100000000010101010010001000100010000000000000000010111011101110110000000000000000";
--X60Y8, nonlinear_LMDPL
constant Tile_X60Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000010101011010101001010101010101010101010100000000101010101100110011001100000000000000000001010101010101010000000000000000";
--X61Y8, linear_LMDPL
constant Tile_X61Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000010101010010001000100010000000000010101010000000000000000001000100010001011011101110111010000000000000000";
--X62Y8, linear_LMDPL
constant Tile_X62Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X63Y8, nonlinear_LMDPL
constant Tile_X63Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010010101011010101000000000101010100000000000000000000000000000000000000000000000001010101010101010010101010101010100000000000000001000100010001000000000000000000001010101010101010000000000000000";
--X64Y8, linear_LMDPL
constant Tile_X64Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X65Y8, linear_LMDPL
constant Tile_X65Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000101010100101010110101010101010100000000000000000111111110000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X66Y8, nonlinear_LMDPL
constant Tile_X66Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111101010101101010100000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111011101110111000000000000000000011001100110011";
--X67Y8, linear_LMDPL
constant Tile_X67Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001111111111111111";
--X68Y8, linear_LMDPL
constant Tile_X68Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X69Y8, nonlinear_LMDPL
constant Tile_X69Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X70Y8, linear_LMDPL
constant Tile_X70Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101011111111100000000101010100000000000000000000000001010101010101010101010100000000001010101000000000000000000000000101010101010101000000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X71Y8, linear_LMDPL
constant Tile_X71Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X72Y8, nonlinear_LMDPL
constant Tile_X72Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X73Y8, linear_LMDPL
constant Tile_X73Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X74Y8, linear_LMDPL
constant Tile_X74Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X75Y8, nonlinear_LMDPL
constant Tile_X75Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000111111110101010100000000010101010101010100000000000000001001100110011001000000000000000011001100110011000000000000000000";
--X76Y8, linear_LMDPL
constant Tile_X76Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X77Y8, linear_LMDPL
constant Tile_X77Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111011101110111010000000000000000";
--X78Y8, ctrl_to_sec
constant Tile_X78Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y8, combined_WDDL
constant Tile_X79Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y8, combined_WDDL
constant Tile_X80Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y8, ctrl_IO
constant Tile_X81Y8_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y9, W_IO_custom
constant Tile_X0Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y9, linear_LMDPL
constant Tile_X1Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X2Y9, linear_LMDPL
constant Tile_X2Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000001010101000000000010101010101010100000000000000001001100110011001000000000000000001000100010001000000000000000000";
--X3Y9, nonlinear_LMDPL
constant Tile_X3Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000111111110000000000000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X4Y9, linear_LMDPL
constant Tile_X4Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001000100010001000000000000000000000010001000100010000000000000000";
--X5Y9, linear_LMDPL
constant Tile_X5Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000011001100110011000110011001100110000000000000000";
--X6Y9, nonlinear_LMDPL
constant Tile_X6Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000010101010110011001100110000000000000000000000000000000000100010001000100";
--X7Y9, linear_LMDPL
constant Tile_X7Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010101010000000010101010111111110000000000000000000000001010101000000000010101010101010100000000000000000001000100010001000000000000000001000100010001000000000000000000";
--X8Y9, linear_LMDPL
constant Tile_X8Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X9Y9, nonlinear_LMDPL
constant Tile_X9Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000010101010000000011111111010101010000000000000000000000001010101000000000000000000000000000000000000000000101010111111111000000001010101000000000010101010101010100000000000000001011101110111011000000000000000000100010001000100000000000000000";
--X10Y9, linear_LMDPL
constant Tile_X10Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000101010100000000000000000000000011111111000000001010101010101010000000000000000000000000000000000101010101010101000000000000000000000000010001000100010000000000010101010000000000000000101110111011101100110011001100110000000000000000";
--X11Y9, linear_LMDPL
constant Tile_X11Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000110011001100110";
--X12Y9, nonlinear_LMDPL
constant Tile_X12Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X13Y9, linear_LMDPL
constant Tile_X13Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001111111111111111";
--X14Y9, linear_LMDPL
constant Tile_X14Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000010101010101010100000000010101010101010100000000010101010101010100000000000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X15Y9, nonlinear_LMDPL
constant Tile_X15Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010011001100110010000000000000000";
--X16Y9, linear_LMDPL
constant Tile_X16Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101010101000000000101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X17Y9, linear_LMDPL
constant Tile_X17Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000101010100000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000010101010111111110000000000000000000100010001000101010101000000001010101010101010000000000000000000000000000000001010101010101010";
--X18Y9, nonlinear_LMDPL
constant Tile_X18Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000101010100000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y9, linear_LMDPL
constant Tile_X19Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000011111111000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X20Y9, linear_LMDPL
constant Tile_X20Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000100010001000100010111011101110110000000000000000";
--X21Y9, nonlinear_LMDPL
constant Tile_X21Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000010101010101010100000000000000001001100110011001000000000000000001000100010001000000000000000000";
--X22Y9, linear_LMDPL
constant Tile_X22Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000000000001010101101010100000000000000000000000000000000000000000101010100101010100000000000000001010101000000000111111110000000010101010010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X23Y9, linear_LMDPL
constant Tile_X23Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001111111111111111";
--X24Y9, nonlinear_LMDPL
constant Tile_X24Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000101010100000000000000000000000001010101000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X25Y9, linear_LMDPL
constant Tile_X25Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010110101010101010101111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X26Y9, linear_LMDPL
constant Tile_X26Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000010101010010001000100010000000000000000000000000000000000110011001100110010111011101110110000000000000000";
--X27Y9, nonlinear_LMDPL
constant Tile_X27Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101011111111101010101010101010101010000000000000000000000000000000000101010101010101000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X28Y9, linear_LMDPL
constant Tile_X28Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000111111111010101000000000000000000000000000000000000000000101010100000000000000001010101010101010000000001010101001010101000000001010101000000000010101010101010110101010000000000011001100110011000000000000000000100010001000100000000000000000";
--X29Y9, linear_LMDPL
constant Tile_X29Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010101010101000000000000000000000000000000000000000000000000101010101111111100000000101010100000000000000000000000001010101010101010010101010000000001010101101010100000000000000000111111110000000010101010010101010101010100000000101010100010001000100010000000000000000011011101110111010000000000000000";
--X30Y9, nonlinear_LMDPL
constant Tile_X30Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010010111011101110110000000000000000";
--X31Y9, linear_LMDPL
constant Tile_X31Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001011101110111011";
--X32Y9, linear_LMDPL
constant Tile_X32Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101010101010101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X33Y9, nonlinear_LMDPL
constant Tile_X33Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101001010101000000000000000010101010000000000101010100000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X34Y9, linear_LMDPL
constant Tile_X34Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000110111011101110110101010101010100000000000000000";
--X35Y9, linear_LMDPL
constant Tile_X35Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010010101010000000001010101000000000000000000000000000000000000000000000000100010001000100000000000000000000010001000100010";
--X36Y9, nonlinear_LMDPL
constant Tile_X36Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000011001100110011";
--X37Y9, linear_LMDPL
constant Tile_X37Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000001010101000000000101010100000000000000000000000001010101000000000101010100101010100000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X38Y9, linear_LMDPL
constant Tile_X38Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000000000000101010100000000000000001010101000000000010001000100010000000000000000000000000000000000110011001100110010001000100010000000000000000000";
--X39Y9, nonlinear_LMDPL
constant Tile_X39Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y9, linear_LMDPL
constant Tile_X40Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010000000001111111100000000010101010101010100000000000000001100110011001100000000000000000001010101010101010000000000000000";
--X41Y9, linear_LMDPL
constant Tile_X41Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010111111111000000000101010100000000101010100000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X42Y9, nonlinear_LMDPL
constant Tile_X42Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000001111111100000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000000000000000000000000000000000000";
--X43Y9, linear_LMDPL
constant Tile_X43Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000001111111100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X44Y9, linear_LMDPL
constant Tile_X44Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101011111111000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000101010101010101010101010101010100000000000000000";
--X45Y9, nonlinear_LMDPL
constant Tile_X45Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010100000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101101010100000000010101010101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X46Y9, linear_LMDPL
constant Tile_X46Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000001010101000000000010101010000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X47Y9, linear_LMDPL
constant Tile_X47Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100101010100000000000000000000000000000000101010100000000011111111010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X48Y9, nonlinear_LMDPL
constant Tile_X48Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000110011001100110";
--X49Y9, linear_LMDPL
constant Tile_X49Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000101010100101010111111111000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X50Y9, linear_LMDPL
constant Tile_X50Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001111111100000000000000000101010111111111000000000000000000000000000000001010101000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X51Y9, nonlinear_LMDPL
constant Tile_X51Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000111111110000000000000000010001000100010000000000010101010000000000000000100110011001100101000100010001000000000000000000";
--X52Y9, linear_LMDPL
constant Tile_X52Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111110101010101010100000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X53Y9, linear_LMDPL
constant Tile_X53Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000111111110000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X54Y9, nonlinear_LMDPL
constant Tile_X54Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X55Y9, linear_LMDPL
constant Tile_X55Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X56Y9, linear_LMDPL
constant Tile_X56Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010111111110000000001010101000000001010101000000000101010100000000000000000000000000101010100000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X57Y9, nonlinear_LMDPL
constant Tile_X57Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001100110011001100000000000000001100110011001100";
--X58Y9, linear_LMDPL
constant Tile_X58Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000110111011101110100000000000000000000000000000000";
--X59Y9, linear_LMDPL
constant Tile_X59Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101011111111010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X60Y9, nonlinear_LMDPL
constant Tile_X60Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000101010100101010100000000000000000000000010101010101010101010101001010101000000000000000011111111000000000000000000000000010001000100010000000000000000001001100110011001";
--X61Y9, linear_LMDPL
constant Tile_X61Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000101010111111111000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000011001100110011";
--X62Y9, linear_LMDPL
constant Tile_X62Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X63Y9, nonlinear_LMDPL
constant Tile_X63Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000010101010000000000000000000000000101010100000000111111110000000010101010010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X64Y9, linear_LMDPL
constant Tile_X64Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X65Y9, linear_LMDPL
constant Tile_X65Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010111111111101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000100010001000100";
--X66Y9, nonlinear_LMDPL
constant Tile_X66Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X67Y9, linear_LMDPL
constant Tile_X67Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X68Y9, linear_LMDPL
constant Tile_X68Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010000000000000000011111111000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X69Y9, nonlinear_LMDPL
constant Tile_X69Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X70Y9, linear_LMDPL
constant Tile_X70Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000001010101101010100000000011111111000000000000000000000000101010100101010101010101000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X71Y9, linear_LMDPL
constant Tile_X71Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110101010100000000000100010001000100000000010101010100010001000100000000000000000000000000000000001100110011001100";
--X72Y9, nonlinear_LMDPL
constant Tile_X72Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X73Y9, linear_LMDPL
constant Tile_X73Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000110011001100110001010101010101010000000000000000";
--X74Y9, linear_LMDPL
constant Tile_X74Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101101010100000000000000000000000000000000010101010000000000000000000000000010101011111111100000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X75Y9, nonlinear_LMDPL
constant Tile_X75Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000000100010001000110111011101110110000000000000000";
--X76Y9, linear_LMDPL
constant Tile_X76Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000001111111100000000010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X77Y9, linear_LMDPL
constant Tile_X77Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000010101010000000000000000011001100110011001110111011101110000000000000000";
--X78Y9, ctrl_to_sec
constant Tile_X78Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y9, combined_WDDL
constant Tile_X79Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000";
--X80Y9, combined_WDDL
constant Tile_X80Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000011110000000011110000000000000000101000000000000000000001000100001010000000000000000000000000111011101110111000000000";
--X81Y9, ctrl_IO
constant Tile_X81Y9_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y10, W_IO_custom
constant Tile_X0Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000";
--X1Y10, linear_LMDPL
constant Tile_X1Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X2Y10, linear_LMDPL
constant Tile_X2Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000001010101000000001010101000000000000000000000000010101010000000000000000000000000110011001100110000000000000000000100010001000100";
--X3Y10, nonlinear_LMDPL
constant Tile_X3Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000010101010000000011111111000000000000000000000000101010100000000000000000010101010101010100000000101010100001000100010001000000000000000000110011001100110000000000000000";
--X4Y10, linear_LMDPL
constant Tile_X4Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000011111111000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X5Y10, linear_LMDPL
constant Tile_X5Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X6Y10, nonlinear_LMDPL
constant Tile_X6Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001110111011101110000000000000000001100110011001100000000000000000";
--X7Y10, linear_LMDPL
constant Tile_X7Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101011111111100000000101010100000000010101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X8Y10, linear_LMDPL
constant Tile_X8Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000010101010000000000000000000000000101010100000000010101010010101010101010100000000000000001111111111111111000000000000000011001100110011000000000000000000";
--X9Y10, nonlinear_LMDPL
constant Tile_X9Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000001000100010001000100010001000100000000000000000";
--X10Y10, linear_LMDPL
constant Tile_X10Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000101010101111111110101010000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X11Y10, linear_LMDPL
constant Tile_X11Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010101010101010101010000000000000000000000000000000000101010100000000111111110000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000101010101010101";
--X12Y10, nonlinear_LMDPL
constant Tile_X12Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X13Y10, linear_LMDPL
constant Tile_X13Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X14Y10, linear_LMDPL
constant Tile_X14Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000010101010101010100000000010101010000000000000000000000000101010101010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X15Y10, nonlinear_LMDPL
constant Tile_X15Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000100010001000100000000101010101001100110011001000000000000000000000000000000001100110011001100";
--X16Y10, linear_LMDPL
constant Tile_X16Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000010101011010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000011001100110011";
--X17Y10, linear_LMDPL
constant Tile_X17Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000111111111010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X18Y10, nonlinear_LMDPL
constant Tile_X18Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010";
--X19Y10, linear_LMDPL
constant Tile_X19Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100101010111111111000000000000000010101010101010100000000010101010010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X20Y10, linear_LMDPL
constant Tile_X20Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X21Y10, nonlinear_LMDPL
constant Tile_X21Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000111111110000000010101010010101010101010100000000101010101101110111011101000000000000000011001100110011000000000000000000";
--X22Y10, linear_LMDPL
constant Tile_X22Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110001010101010101010000000000000000";
--X23Y10, linear_LMDPL
constant Tile_X23Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000010101010101010100000000000000000010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X24Y10, nonlinear_LMDPL
constant Tile_X24Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111111111111000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X25Y10, linear_LMDPL
constant Tile_X25Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000101010100101010110101010010101010101010100000000000000001100110011001100000000000000000010111011101110110000000000000000";
--X26Y10, linear_LMDPL
constant Tile_X26Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X27Y10, nonlinear_LMDPL
constant Tile_X27Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000001010101101010100000000000000000000000001010101000000000010101011010101010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010010111011101110110000000000000000";
--X28Y10, linear_LMDPL
constant Tile_X28Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X29Y10, linear_LMDPL
constant Tile_X29Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000101010101010101011111111101010100000000001010101000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001011101110111011";
--X30Y10, nonlinear_LMDPL
constant Tile_X30Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X31Y10, linear_LMDPL
constant Tile_X31Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101011111111101010100000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X32Y10, linear_LMDPL
constant Tile_X32Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101011111111101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X33Y10, nonlinear_LMDPL
constant Tile_X33Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100101010110101010000000000000000000000000000000000000000010101010000100010001000100000000101010101011101110111011000000000000000000000000000000000011001100110011";
--X34Y10, linear_LMDPL
constant Tile_X34Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000101010100000000000000000000000000000000101010100000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000101010101010101000000000000000000000000000000001100110011001100";
--X35Y10, linear_LMDPL
constant Tile_X35Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010110101010000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X36Y10, nonlinear_LMDPL
constant Tile_X36Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000001010101000000000101010100000000000000000000100010001000100000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X37Y10, linear_LMDPL
constant Tile_X37Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010101010101000000000000000000000000000000000000000000101010101010101101010100000000001010101101010100000000000000000101010100000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000011101110111011100000000000000001100110011001100";
--X38Y10, linear_LMDPL
constant Tile_X38Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X39Y10, nonlinear_LMDPL
constant Tile_X39Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010011001100110010000000000000000";
--X40Y10, linear_LMDPL
constant Tile_X40Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001110111011101110000000000000000";
--X41Y10, linear_LMDPL
constant Tile_X41Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X42Y10, nonlinear_LMDPL
constant Tile_X42Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000000000001010101011111111000000001010101000000000000000000000000000000000010101010101010100000000101010100001000100010001000000000000000001000100010001000000000000000000";
--X43Y10, linear_LMDPL
constant Tile_X43Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101111111100000000101010100000000000000000000000001010101010101010000000000000000010101010000000000101010111111111010101010101010100000000000000000111011101110111000000000000000010111011101110110000000000000000";
--X44Y10, linear_LMDPL
constant Tile_X44Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010101010101010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X45Y10, nonlinear_LMDPL
constant Tile_X45Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000010001000100010000010001000100010000000000000000";
--X46Y10, linear_LMDPL
constant Tile_X46Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000010101010000000001010101000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000010101010101010100100010001000100000000000000000";
--X47Y10, linear_LMDPL
constant Tile_X47Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X48Y10, nonlinear_LMDPL
constant Tile_X48Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000101010101010101010011001100110010000000000000000";
--X49Y10, linear_LMDPL
constant Tile_X49Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101011010101000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101011111111010101010101010100000000000000000100010001000100000000000000000001110111011101110000000000000000";
--X50Y10, linear_LMDPL
constant Tile_X50Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000101010100000000010101010101010100000000101010101011101110111011000000000000000010001000100010000000000000000000";
--X51Y10, nonlinear_LMDPL
constant Tile_X51Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X52Y10, linear_LMDPL
constant Tile_X52Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X53Y10, linear_LMDPL
constant Tile_X53Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110111011101110100000000000000000000000000000000";
--X54Y10, nonlinear_LMDPL
constant Tile_X54Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000001010101000000000101010100000000101010101010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000100010001000100";
--X55Y10, linear_LMDPL
constant Tile_X55Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001000100010001000";
--X56Y10, linear_LMDPL
constant Tile_X56Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000101010100000000000000000101010101010101000000000000000000100010001000100";
--X57Y10, nonlinear_LMDPL
constant Tile_X57Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000101010100000000000100010001000100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X58Y10, linear_LMDPL
constant Tile_X58Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000001010101001010101101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X59Y10, linear_LMDPL
constant Tile_X59Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000101010101101110111011101000000000000000001010101010101010000000000000000";
--X60Y10, nonlinear_LMDPL
constant Tile_X60Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000001010101000000000000000000000000101010100000000000000000000000000101010111111111000000000000000010101010010101010101010100000000101010101001100110011001000000000000000010111011101110110000000000000000";
--X61Y10, linear_LMDPL
constant Tile_X61Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000101010100100010001000100000000000000000000000000000000000011001100110011";
--X62Y10, linear_LMDPL
constant Tile_X62Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101011010101000000000000000000000000010101010000000001010101000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X63Y10, nonlinear_LMDPL
constant Tile_X63Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X64Y10, linear_LMDPL
constant Tile_X64Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111111111111100000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111111111111111100000000000000000000000000000000";
--X65Y10, linear_LMDPL
constant Tile_X65Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001101110111011101";
--X66Y10, nonlinear_LMDPL
constant Tile_X66Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000011101110111011100000000000000000";
--X67Y10, linear_LMDPL
constant Tile_X67Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000100010001000100";
--X68Y10, linear_LMDPL
constant Tile_X68Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000001010101010101010000000000000000011111111000000000000000000000000111111110101010100000000010101010101010100000000000000000111011101110111000000000000000010001000100010000000000000000000";
--X69Y10, nonlinear_LMDPL
constant Tile_X69Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111000000000000000000000000010101010000000010101010010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X70Y10, linear_LMDPL
constant Tile_X70Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000111111111010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000001000100010001";
--X71Y10, linear_LMDPL
constant Tile_X71Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010101010100000000000000000000000001111111100000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X72Y10, nonlinear_LMDPL
constant Tile_X72Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X73Y10, linear_LMDPL
constant Tile_X73Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101011111111000000000000000000000000010101010000000000000000010001000100010000000000111111110000000000000000000100010001000100110011001100110000000000000000";
--X74Y10, linear_LMDPL
constant Tile_X74Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001111111101010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000001010101010101010000000000000000";
--X75Y10, nonlinear_LMDPL
constant Tile_X75Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000100010001000100000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X76Y10, linear_LMDPL
constant Tile_X76Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X77Y10, linear_LMDPL
constant Tile_X77Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000010101010000000000000000000000000000000011111111111111110000000000000000";
--X78Y10, ctrl_to_sec
constant Tile_X78Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y10, combined_WDDL
constant Tile_X79Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y10, combined_WDDL
constant Tile_X80Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y10, ctrl_IO
constant Tile_X81Y10_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y11, W_IO_custom
constant Tile_X0Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y11, linear_LMDPL
constant Tile_X1Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011101110111011100000000000000000000000000000000";
--X2Y11, linear_LMDPL
constant Tile_X2Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000111111111111111101000100010001000000000000000000";
--X3Y11, nonlinear_LMDPL
constant Tile_X3Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001111111100000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X4Y11, linear_LMDPL
constant Tile_X4Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001100110011001100000000000000000";
--X5Y11, linear_LMDPL
constant Tile_X5Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000001010101010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X6Y11, nonlinear_LMDPL
constant Tile_X6Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000111111110000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001001100110011001";
--X7Y11, linear_LMDPL
constant Tile_X7Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000001010101011111111010101010101010100000000000000000110011001100110000000000000000001010101010101010000000000000000";
--X8Y11, linear_LMDPL
constant Tile_X8Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000001100110011001110101010101010100000000000000000";
--X9Y11, nonlinear_LMDPL
constant Tile_X9Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000111111110000000000000000000000000000000011111111000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001100110011001100";
--X10Y11, linear_LMDPL
constant Tile_X10Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000010101010000000001010101000000000010101010000000000000000111111110000000000000000000000000000000001010101010101010101010100000000000000000011001100110011000000000000000011011101110111010000000000000000";
--X11Y11, linear_LMDPL
constant Tile_X11Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000011001100110011000000000000000011101110111011100000000000000000";
--X12Y11, nonlinear_LMDPL
constant Tile_X12Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000001010101000000001111111100000000101010101010101000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X13Y11, linear_LMDPL
constant Tile_X13Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X14Y11, linear_LMDPL
constant Tile_X14Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100000000010101010000000000000000000000000101010101010101000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001011101110111011";
--X15Y11, nonlinear_LMDPL
constant Tile_X15Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000001010101011111111000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X16Y11, linear_LMDPL
constant Tile_X16Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X17Y11, linear_LMDPL
constant Tile_X17Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X18Y11, nonlinear_LMDPL
constant Tile_X18Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X19Y11, linear_LMDPL
constant Tile_X19Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000101010101010101000000000000000000000000101010101010101000000000010101010000000000000000000000000000000000000000000000001111111110101010010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X20Y11, linear_LMDPL
constant Tile_X20Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000001010101000000000101010101010101010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000010101010010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X21Y11, nonlinear_LMDPL
constant Tile_X21Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000010101010010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X22Y11, linear_LMDPL
constant Tile_X22Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000001010101000000000000000000000000011111111010101010101010111111111000000000100010001000100000000000000000001110111011101110000000000000000";
--X23Y11, linear_LMDPL
constant Tile_X23Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010100000000011111111010101010101010100000000000000000101010101010101000000000000000010001000100010000000000000000000";
--X24Y11, nonlinear_LMDPL
constant Tile_X24Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101011010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X25Y11, linear_LMDPL
constant Tile_X25Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000010001000100010010111011101110110000000000000000";
--X26Y11, linear_LMDPL
constant Tile_X26Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X27Y11, nonlinear_LMDPL
constant Tile_X27Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010010101010000000000000000000000001010101000000000000000000101010110101010000000000000000000000000010101010000000010101010010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X28Y11, linear_LMDPL
constant Tile_X28Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000001111111100000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010000000001111111110101010000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X29Y11, linear_LMDPL
constant Tile_X29Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000110111011101110100000000000000001111111111111111";
--X30Y11, nonlinear_LMDPL
constant Tile_X30Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000101010100000000101010100101010111111111000000000101010110101010000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X31Y11, linear_LMDPL
constant Tile_X31Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101011111111101010100101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001000100010001000";
--X32Y11, linear_LMDPL
constant Tile_X32Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010101010100000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000101010101010101011111111101010100101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000001011101110111011";
--X33Y11, nonlinear_LMDPL
constant Tile_X33Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101010101010000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000000001000100010001";
--X34Y11, linear_LMDPL
constant Tile_X34Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000111111111111111110101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001010101010101010000000000000000";
--X35Y11, linear_LMDPL
constant Tile_X35Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010111111110000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X36Y11, nonlinear_LMDPL
constant Tile_X36Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000001010101010101010";
--X37Y11, linear_LMDPL
constant Tile_X37Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X38Y11, linear_LMDPL
constant Tile_X38Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000101010100101010100000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X39Y11, nonlinear_LMDPL
constant Tile_X39Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X40Y11, linear_LMDPL
constant Tile_X40Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000101010101010101000000000000000000100010001000100";
--X41Y11, linear_LMDPL
constant Tile_X41Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000010101010010101010101010111111111000000000000000000000000000000000000000001000100010001000000000000000000";
--X42Y11, nonlinear_LMDPL
constant Tile_X42Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010101010000000010101010000000000000000000000000000000000000000011111111010001000100010000000000101010100000000000000000100010001000100010011001100110010000000000000000";
--X43Y11, linear_LMDPL
constant Tile_X43Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000101010110101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001011101110111011000000000000000000100010001000100000000000000000";
--X44Y11, linear_LMDPL
constant Tile_X44Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101011011101110111010000000000000000";
--X45Y11, nonlinear_LMDPL
constant Tile_X45Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000000100010001000100100010001000100000000000000000";
--X46Y11, linear_LMDPL
constant Tile_X46Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000001010101000000001010101010101010000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X47Y11, linear_LMDPL
constant Tile_X47Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000011101110111011100000000000000000010001000100010";
--X48Y11, nonlinear_LMDPL
constant Tile_X48Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110000000000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000100010001000100";
--X49Y11, linear_LMDPL
constant Tile_X49Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000111111110000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000101010101000100010001000000000000000000000000000000000000011001100110011";
--X50Y11, linear_LMDPL
constant Tile_X50Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001111111101010101101010100000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X51Y11, nonlinear_LMDPL
constant Tile_X51Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000101010100000000000000001010101000000000010101010000000000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000110011001100110";
--X52Y11, linear_LMDPL
constant Tile_X52Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010101010100000000000000000101010101010101000000000000000000000000001010101000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X53Y11, linear_LMDPL
constant Tile_X53Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000101010101111111100000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000";
--X54Y11, nonlinear_LMDPL
constant Tile_X54Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100000000000000000111111110000000000000000010101010000000000000000000000000000000000000000101010101010101000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000010001000100010";
--X55Y11, linear_LMDPL
constant Tile_X55Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X56Y11, linear_LMDPL
constant Tile_X56Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000010101010000000001010101001010101101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X57Y11, nonlinear_LMDPL
constant Tile_X57Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000001010101111111110000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001000100010001000";
--X58Y11, linear_LMDPL
constant Tile_X58Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000111111110101010100000000000000000000000010101010000000000101010100000000000000000000000001010101000000000000000000000000101010100000000000000000010001000100010000000000000000001100110011001100";
--X59Y11, linear_LMDPL
constant Tile_X59Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X60Y11, nonlinear_LMDPL
constant Tile_X60Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010101010010101010101010100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X61Y11, linear_LMDPL
constant Tile_X61Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010011111111000000000000000000000000001000100010001010001000100010000000000000000000";
--X62Y11, linear_LMDPL
constant Tile_X62Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000001111111110101010000000000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X63Y11, nonlinear_LMDPL
constant Tile_X63Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X64Y11, linear_LMDPL
constant Tile_X64Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000011111111101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X65Y11, linear_LMDPL
constant Tile_X65Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001111111111111111";
--X66Y11, nonlinear_LMDPL
constant Tile_X66Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X67Y11, linear_LMDPL
constant Tile_X67Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X68Y11, linear_LMDPL
constant Tile_X68Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010101010101010101010000000000000000011111111000000000000000000000000101010100101010110101010010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X69Y11, nonlinear_LMDPL
constant Tile_X69Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000100010001000100000000010101011100110011001100000000000000000000000000000000000000000000000000";
--X70Y11, linear_LMDPL
constant Tile_X70Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000000000000011111111000000001010101010101010010001000100010011111111000000000000000000000000001000100010001011001100110011000000000000000000";
--X71Y11, linear_LMDPL
constant Tile_X71Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000000100010001000100000000000000000010001000100010";
--X72Y11, nonlinear_LMDPL
constant Tile_X72Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000010101010010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X73Y11, linear_LMDPL
constant Tile_X73Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000101010100101010101010101000000000000000010011001100110010000000000000000";
--X74Y11, linear_LMDPL
constant Tile_X74Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000010101010101010100000000010101011000100010001000000000000000000000000000000000000000000000000000";
--X75Y11, nonlinear_LMDPL
constant Tile_X75Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000010101010011001100110011000000000000000000000000000000000001000100010001";
--X76Y11, linear_LMDPL
constant Tile_X76Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000001000100010001000000000000000001011101110111011";
--X77Y11, linear_LMDPL
constant Tile_X77Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000010101010000000000000000001100110011001110101010101010100000000000000000";
--X78Y11, ctrl_to_sec
constant Tile_X78Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y11, combined_WDDL
constant Tile_X79Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y11, combined_WDDL
constant Tile_X80Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y11, ctrl_IO
constant Tile_X81Y11_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y12, W_IO_custom
constant Tile_X0Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000";
--X1Y12, linear_LMDPL
constant Tile_X1Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001001100110011001";
--X2Y12, linear_LMDPL
constant Tile_X2Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X3Y12, nonlinear_LMDPL
constant Tile_X3Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000001000100010001";
--X4Y12, linear_LMDPL
constant Tile_X4Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000001010101000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X5Y12, linear_LMDPL
constant Tile_X5Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X6Y12, nonlinear_LMDPL
constant Tile_X6Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X7Y12, linear_LMDPL
constant Tile_X7Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X8Y12, linear_LMDPL
constant Tile_X8Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110000000000000000010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X9Y12, nonlinear_LMDPL
constant Tile_X9Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101010101010000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X10Y12, linear_LMDPL
constant Tile_X10Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010101010100000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000011011101110111010000000000000000";
--X11Y12, linear_LMDPL
constant Tile_X11Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101011010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001010101010101010";
--X12Y12, nonlinear_LMDPL
constant Tile_X12Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X13Y12, linear_LMDPL
constant Tile_X13Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000001111111100000000010001000100010000000000000000000000000000000000101110111011101110111011101110110000000000000000";
--X14Y12, linear_LMDPL
constant Tile_X14Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010101111111110101010101010100000000001010101101010101010101000000000010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X15Y12, nonlinear_LMDPL
constant Tile_X15Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000100010001000100010011001100110010000000000000000";
--X16Y12, linear_LMDPL
constant Tile_X16Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000010101011010101010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X17Y12, linear_LMDPL
constant Tile_X17Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000100010001000100000000000000001111111111111111000000000000000000000000000000000101010101010101";
--X18Y12, nonlinear_LMDPL
constant Tile_X18Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y12, linear_LMDPL
constant Tile_X19Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010101010100000000010101010000100010001000100000000000000001011101110111011000000000000000000000000000000000001000100010001";
--X20Y12, linear_LMDPL
constant Tile_X20Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000011111111000000000000000000000000101010100000000010101010010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X21Y12, nonlinear_LMDPL
constant Tile_X21Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000101010100001000100010001000000000000000010101010101010100000000000000000";
--X22Y12, linear_LMDPL
constant Tile_X22Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110010101010101010100000000000000000";
--X23Y12, linear_LMDPL
constant Tile_X23Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000001010101000000000000000000101010100000000010101010000000010101010101010100000000000000000010001000100010000000000000000000000000000000000110111011101110110101010101010100000000000000000";
--X24Y12, nonlinear_LMDPL
constant Tile_X24Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X25Y12, linear_LMDPL
constant Tile_X25Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X26Y12, linear_LMDPL
constant Tile_X26Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X27Y12, nonlinear_LMDPL
constant Tile_X27Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000010101010000000000000000000000000000000000101010100000000000000001010101010101010000000000000000000000000111111110000000010101010010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X28Y12, linear_LMDPL
constant Tile_X28Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000110101010000000000000000000000000000000000000000000000000000000001010101010101010";
--X29Y12, linear_LMDPL
constant Tile_X29Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000101010100000000000000000101010101111111100000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X30Y12, nonlinear_LMDPL
constant Tile_X30Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X31Y12, linear_LMDPL
constant Tile_X31Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000001010101101010100000000000000000010101011010101000000000101010100000000000000000111111110000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X32Y12, linear_LMDPL
constant Tile_X32Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000111111111010101010101010101010101010101000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110100100010001000100000000000000000";
--X33Y12, nonlinear_LMDPL
constant Tile_X33Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000101010100000000000000000000000001010101000000000101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X34Y12, linear_LMDPL
constant Tile_X34Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X35Y12, linear_LMDPL
constant Tile_X35Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000001010101000000000101010100000000000000000000000000000000000000000010101010000000000000000100010001000100000000000000000001010101010101010";
--X36Y12, nonlinear_LMDPL
constant Tile_X36Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000011001100110011";
--X37Y12, linear_LMDPL
constant Tile_X37Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010000000000000000000000001010101000000000000000000000000011111111000100010001000100000000000000001100110011001100000000000000000000000000000000001111111111111111";
--X38Y12, linear_LMDPL
constant Tile_X38Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100101010100000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000011001100110011011001100110011000000000000000000";
--X39Y12, nonlinear_LMDPL
constant Tile_X39Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000101010100000000101010100000000000000000010001000100010000000000101010100000000000000000100110011001100110101010101010100000000000000000";
--X40Y12, linear_LMDPL
constant Tile_X40Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000010101010000000000000000000000000000000001010101000000000000000000000000101010100000000000000000101010100000000000000000101010100101010100000000000000000000000010101010000000000000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X41Y12, linear_LMDPL
constant Tile_X41Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X42Y12, nonlinear_LMDPL
constant Tile_X42Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000101010100000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001000100010001000";
--X43Y12, linear_LMDPL
constant Tile_X43Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010110101010101010100000000000000000010101010000000000000000101010100000000000000000000000000000000001010101000000001010101000000000010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X44Y12, linear_LMDPL
constant Tile_X44Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010101011010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001010001000100010000000000000000000";
--X45Y12, nonlinear_LMDPL
constant Tile_X45Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010101010101000000000000000000000000000000000000000011111111010101010101010100000000101010101100110011001100000000000000000010101010101010100000000000000000";
--X46Y12, linear_LMDPL
constant Tile_X46Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000001010101000000000000000000000000101010101111111100000000000000001010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X47Y12, linear_LMDPL
constant Tile_X47Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101001010101000000000000000000000000000000000000000011111111010101010000000011111111000000000000000000000000101010100000000001010101010101010101010100000000000000001100110011001100000000000000000001010101010101010000000000000000";
--X48Y12, nonlinear_LMDPL
constant Tile_X48Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000001000100010001";
--X49Y12, linear_LMDPL
constant Tile_X49Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X50Y12, linear_LMDPL
constant Tile_X50Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000101010100000000000000000101010100000000001010101000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010101010101010100000000101010100101010101010101000000000000000010001000100010000000000000000000";
--X51Y12, nonlinear_LMDPL
constant Tile_X51Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101000000000000000001010101000000000111111110000000010101010010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X52Y12, linear_LMDPL
constant Tile_X52Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101010101010101010100101010111111111000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X53Y12, linear_LMDPL
constant Tile_X53Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000010101010000000000000000000000000101010100000000000000000101010100101010100000000101010100000000000000000000000000000000010101010010101010000000010101010010101010101010100000000101010100101010101010101000000000000000000000000000000000000000000000000";
--X54Y12, nonlinear_LMDPL
constant Tile_X54Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000001111111100000000000000000000000000000000101010100000000000000000101010101010101000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010101010100000000010101011011101110111011000000000000000000000000000000000000000000000000";
--X55Y12, linear_LMDPL
constant Tile_X55Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X56Y12, linear_LMDPL
constant Tile_X56Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X57Y12, nonlinear_LMDPL
constant Tile_X57Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000001111111100000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X58Y12, linear_LMDPL
constant Tile_X58Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000101010110101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X59Y12, linear_LMDPL
constant Tile_X59Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000001010101010101010101010100000000101010101011101110111011000000000000000011001100110011000000000000000000";
--X60Y12, nonlinear_LMDPL
constant Tile_X60Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000101010100000000111111110000000000000000010101010101010100000000101010101111111111111111000000000000000011011101110111010000000000000000";
--X61Y12, linear_LMDPL
constant Tile_X61Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X62Y12, linear_LMDPL
constant Tile_X62Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X63Y12, nonlinear_LMDPL
constant Tile_X63Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111101010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X64Y12, linear_LMDPL
constant Tile_X64Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000101010100000000000000000111111110000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000110011001100110011001100110011000000000000000000";
--X65Y12, linear_LMDPL
constant Tile_X65Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010110101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X66Y12, nonlinear_LMDPL
constant Tile_X66Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001010101000000001111111110101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000110011001100110000000000000000000100010001000100";
--X67Y12, linear_LMDPL
constant Tile_X67Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X68Y12, linear_LMDPL
constant Tile_X68Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000101010111111111000000001010101010101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X69Y12, nonlinear_LMDPL
constant Tile_X69Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000101010110101010010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X70Y12, linear_LMDPL
constant Tile_X70Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101111111110101010000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X71Y12, linear_LMDPL
constant Tile_X71Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000010101010000000000000000101010101010101001000100010001000000000000000000";
--X72Y12, nonlinear_LMDPL
constant Tile_X72Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000010101011000100010001000000000000000000010101010101010100000000000000000";
--X73Y12, linear_LMDPL
constant Tile_X73Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101011110111011101110000000000000000000100010001000100000000000000000";
--X74Y12, linear_LMDPL
constant Tile_X74Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001000100010001000";
--X75Y12, nonlinear_LMDPL
constant Tile_X75Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000101010101000100010001000000000000000000010011001100110010000000000000000";
--X76Y12, linear_LMDPL
constant Tile_X76Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X77Y12, linear_LMDPL
constant Tile_X77Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000001100110011001100000000000000000000000000000000";
--X78Y12, ctrl_to_sec
constant Tile_X78Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y12, combined_WDDL
constant Tile_X79Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y12, combined_WDDL
constant Tile_X80Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y12, ctrl_IO
constant Tile_X81Y12_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y13, W_IO_custom
constant Tile_X0Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001111111110000000000010101010000000000000000000000000";
--X1Y13, linear_LMDPL
constant Tile_X1Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000111011101110111";
--X2Y13, linear_LMDPL
constant Tile_X2Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X3Y13, nonlinear_LMDPL
constant Tile_X3Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000100010001000100000000000000000";
--X4Y13, linear_LMDPL
constant Tile_X4Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000010101010000000010101010010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X5Y13, linear_LMDPL
constant Tile_X5Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010101111111100000000000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X6Y13, nonlinear_LMDPL
constant Tile_X6Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000100010001000100000010001000100010000000000000000";
--X7Y13, linear_LMDPL
constant Tile_X7Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111010101010101010100000000111111110100010001000100000000000000000011001100110011000000000000000000";
--X8Y13, linear_LMDPL
constant Tile_X8Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X9Y13, nonlinear_LMDPL
constant Tile_X9Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X10Y13, linear_LMDPL
constant Tile_X10Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111010101011010101000000000000000000000000000000000000000001010101001010101010101010101010100000000101010100000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X11Y13, linear_LMDPL
constant Tile_X11Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000100010001000100000000000000000000101010101010101";
--X12Y13, nonlinear_LMDPL
constant Tile_X12Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000001111111100000000010001000100010000000000000000000000000000000000001000100010001000010001000100010000000000000000";
--X13Y13, linear_LMDPL
constant Tile_X13Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X14Y13, linear_LMDPL
constant Tile_X14Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100";
--X15Y13, nonlinear_LMDPL
constant Tile_X15Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000001000100010001";
--X16Y13, linear_LMDPL
constant Tile_X16Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X17Y13, linear_LMDPL
constant Tile_X17Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X18Y13, nonlinear_LMDPL
constant Tile_X18Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000001000100010001000000000000000000001000100010001";
--X19Y13, linear_LMDPL
constant Tile_X19Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X20Y13, linear_LMDPL
constant Tile_X20Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X21Y13, nonlinear_LMDPL
constant Tile_X21Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X22Y13, linear_LMDPL
constant Tile_X22Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000111011101110111000000000000000000000000000000000000000000000000";
--X23Y13, linear_LMDPL
constant Tile_X23Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000001111111100000000000000001010101011111111000000000000000000000000010101010000000000000000010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X24Y13, nonlinear_LMDPL
constant Tile_X24Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X25Y13, linear_LMDPL
constant Tile_X25Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X26Y13, linear_LMDPL
constant Tile_X26Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X27Y13, nonlinear_LMDPL
constant Tile_X27Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X28Y13, linear_LMDPL
constant Tile_X28Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110111011101110111011101110111010000000000000000";
--X29Y13, linear_LMDPL
constant Tile_X29Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001010101010101010";
--X30Y13, nonlinear_LMDPL
constant Tile_X30Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100101010110101010000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y13, linear_LMDPL
constant Tile_X31Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000101010100000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X32Y13, linear_LMDPL
constant Tile_X32Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100101010100000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010101010100000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X33Y13, nonlinear_LMDPL
constant Tile_X33Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000001010101000000000101010100101010100000000000000000000000000000000010101010000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000001100110011001100";
--X34Y13, linear_LMDPL
constant Tile_X34Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X35Y13, linear_LMDPL
constant Tile_X35Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000010101010010101010000000010101010000000000000000000000000101010100000000011111111000100010001000100000000010101011101110111011101000000000000000000000000000000001010101010101010";
--X36Y13, nonlinear_LMDPL
constant Tile_X36Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001000100010001000";
--X37Y13, linear_LMDPL
constant Tile_X37Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X38Y13, linear_LMDPL
constant Tile_X38Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000001010101000000000101010100000000001010101000000000000000000000000000000000000000000000000010101010101010100000000010101010100010001000100000000000000000010111011101110110000000000000000";
--X39Y13, nonlinear_LMDPL
constant Tile_X39Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000101010100000000000000000010101011010101000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000010101010101010100000000000000000001000100010001000000000000000001010101010101010000000000000000";
--X40Y13, linear_LMDPL
constant Tile_X40Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000101010101010101000000000000000001010101000000000000000000101010110101010000000000000000001010101010101010101010100000000000000000101010101010101000000000000000010101010101010100000000000000000";
--X41Y13, linear_LMDPL
constant Tile_X41Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100101010110101010000000000000000001010101101010100000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X42Y13, nonlinear_LMDPL
constant Tile_X42Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010111111110000000000000000101010100000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000001101110111011101";
--X43Y13, linear_LMDPL
constant Tile_X43Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000101010101010101101010100000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000011001100110011000000000000000000011001100110011";
--X44Y13, linear_LMDPL
constant Tile_X44Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X45Y13, nonlinear_LMDPL
constant Tile_X45Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000001010101000000000000000001010101010101010000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X46Y13, linear_LMDPL
constant Tile_X46Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000000000000010101011010101010101010000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X47Y13, linear_LMDPL
constant Tile_X47Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000001111111100000000000000001010101000000000000000000000000001010101000000000000000000000000000000000101010110101010000000000000000000000000000000000000000001010101010101010101010100000000010101011100110011001100000000000000000001110111011101110000000000000000";
--X48Y13, nonlinear_LMDPL
constant Tile_X48Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X49Y13, linear_LMDPL
constant Tile_X49Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010010101010101010100000000101010100000000000000000000000000000000010001000100010000000000000000000";
--X50Y13, linear_LMDPL
constant Tile_X50Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010101010101111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X51Y13, nonlinear_LMDPL
constant Tile_X51Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000001010101000000000000000001010101000000000111111110101010110101010010001000100010000000000010101010000000000000000101010101010101011001100110011000000000000000000";
--X52Y13, linear_LMDPL
constant Tile_X52Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111110101010101010100101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X53Y13, linear_LMDPL
constant Tile_X53Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101011111111101010101010101010000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010100000000000000000111111110101010100000000000000000000000000000000010101010101010110101010000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X54Y13, nonlinear_LMDPL
constant Tile_X54Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000100110011001100100100010001000100000000000000000";
--X55Y13, linear_LMDPL
constant Tile_X55Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000001010101000000000111111110000000000000000101010100000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X56Y13, linear_LMDPL
constant Tile_X56Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X57Y13, nonlinear_LMDPL
constant Tile_X57Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X58Y13, linear_LMDPL
constant Tile_X58Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000111111110000000011111111000000000000000011111111000000000000000010101010010101010101010100000000101010100010001000100010000000000000000000000000000000000000000000000000";
--X59Y13, linear_LMDPL
constant Tile_X59Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000011111111010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X60Y13, nonlinear_LMDPL
constant Tile_X60Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000001010101101010100000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000101010111111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X61Y13, linear_LMDPL
constant Tile_X61Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000001000100010001000000000000000000";
--X62Y13, linear_LMDPL
constant Tile_X62Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111110101010000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X63Y13, nonlinear_LMDPL
constant Tile_X63Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111110101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000010101011010101010101010000000000000000000100010001000100000000000000000";
--X64Y13, linear_LMDPL
constant Tile_X64Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010000000000000000111111110000000000000000101010100000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000100010001000100";
--X65Y13, linear_LMDPL
constant Tile_X65Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001111111111111111101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X66Y13, nonlinear_LMDPL
constant Tile_X66Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X67Y13, linear_LMDPL
constant Tile_X67Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X68Y13, linear_LMDPL
constant Tile_X68Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101010101010000000000101010100000000000000000000000000000000000000000101010111111111010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X69Y13, nonlinear_LMDPL
constant Tile_X69Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000101010101111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000010101011010101010101010000000000000000011001100110011000000000000000000";
--X70Y13, linear_LMDPL
constant Tile_X70Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000101010100000000010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X71Y13, linear_LMDPL
constant Tile_X71Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000111111111010101000000000000000001010101000000000000000000000000010101010000100010001000100000000010101011001100110011001000000000000000000000000000000000010001000100010";
--X72Y13, nonlinear_LMDPL
constant Tile_X72Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X73Y13, linear_LMDPL
constant Tile_X73Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000010001000100010";
--X74Y13, linear_LMDPL
constant Tile_X74Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000101010100000000101010101010101011111111010101010101010100000000101010101100110011001100000000000000000000000000000000000000000000000000";
--X75Y13, nonlinear_LMDPL
constant Tile_X75Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000101010101000100010001000000000000000000001010101010101010000000000000000";
--X76Y13, linear_LMDPL
constant Tile_X76Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000000000000000000010111011101110110000000000000000";
--X77Y13, linear_LMDPL
constant Tile_X77Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010101010100000000101010101000100010001000000000000000000010111011101110110000000000000000";
--X78Y13, ctrl_to_sec
constant Tile_X78Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y13, combined_WDDL
constant Tile_X79Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y13, combined_WDDL
constant Tile_X80Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y13, ctrl_IO
constant Tile_X81Y13_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y14, W_IO_custom
constant Tile_X0Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000100100100101000000000000000010100000000000000000000000000000000";
--X1Y14, linear_LMDPL
constant Tile_X1Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010101111111100000000010001000100010000000000000000000000000000000000010101010101010101000100010001000000000000000000";
--X2Y14, linear_LMDPL
constant Tile_X2Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000001010101000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X3Y14, nonlinear_LMDPL
constant Tile_X3Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000101010101010101000010001000100010000000000000000";
--X4Y14, linear_LMDPL
constant Tile_X4Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X5Y14, linear_LMDPL
constant Tile_X5Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X6Y14, nonlinear_LMDPL
constant Tile_X6Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000000000001010101010101010000000000000000001110111011101110000000000000000";
--X7Y14, linear_LMDPL
constant Tile_X7Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X8Y14, linear_LMDPL
constant Tile_X8Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000111111110000000000000000010001000100010000000000111111110000000000000000001000100010001001010101010101010000000000000000";
--X9Y14, nonlinear_LMDPL
constant Tile_X9Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000010001000100010";
--X10Y14, linear_LMDPL
constant Tile_X10Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X11Y14, linear_LMDPL
constant Tile_X11Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000111011101110111000000000000000000000000000000000000000000000000";
--X12Y14, nonlinear_LMDPL
constant Tile_X12Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001011101110111011";
--X13Y14, linear_LMDPL
constant Tile_X13Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X14Y14, linear_LMDPL
constant Tile_X14Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100000000010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X15Y14, nonlinear_LMDPL
constant Tile_X15Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X16Y14, linear_LMDPL
constant Tile_X16Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X17Y14, linear_LMDPL
constant Tile_X17Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001110111011101110";
--X18Y14, nonlinear_LMDPL
constant Tile_X18Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010011001100110010000000000000000";
--X19Y14, linear_LMDPL
constant Tile_X19Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000011001100110011";
--X20Y14, linear_LMDPL
constant Tile_X20Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X21Y14, nonlinear_LMDPL
constant Tile_X21Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000111011101110111000000000000000000101010101010101";
--X22Y14, linear_LMDPL
constant Tile_X22Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000010101010101010100000000101010101111111111111111000000000000000001000100010001000000000000000000";
--X23Y14, linear_LMDPL
constant Tile_X23Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X24Y14, nonlinear_LMDPL
constant Tile_X24Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000001001100110011001";
--X25Y14, linear_LMDPL
constant Tile_X25Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X26Y14, linear_LMDPL
constant Tile_X26Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X27Y14, nonlinear_LMDPL
constant Tile_X27Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000111111110000000010101010010001000100010000000000010101010000000000000000001100110011001110011001100110010000000000000000";
--X28Y14, linear_LMDPL
constant Tile_X28Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000101010101010101000000000000000011001100110011000000000000000000";
--X29Y14, linear_LMDPL
constant Tile_X29Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000111111110101010100000000111111110000000000000000101010100000000001010101000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X30Y14, nonlinear_LMDPL
constant Tile_X30Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101010101010000000000000000000000000000000001010101000000000101010100101010110101010000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000100010001000100";
--X31Y14, linear_LMDPL
constant Tile_X31Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101111111101010101010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100101010100000000111111110000000010101010101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001101110111011101";
--X32Y14, linear_LMDPL
constant Tile_X32Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X33Y14, nonlinear_LMDPL
constant Tile_X33Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000101010100101010100000000000000000000000000000000000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000100010001000100";
--X34Y14, linear_LMDPL
constant Tile_X34Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000010101010000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X35Y14, linear_LMDPL
constant Tile_X35Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000010101010000000000000000010101010111111110000000010101010000000001010101000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X36Y14, nonlinear_LMDPL
constant Tile_X36Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101111111100000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010100101010100000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000010001000100010";
--X37Y14, linear_LMDPL
constant Tile_X37Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000111011101110111";
--X38Y14, linear_LMDPL
constant Tile_X38Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000011111111000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X39Y14, nonlinear_LMDPL
constant Tile_X39Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000101010100111011101110111000000000000000011001100110011000000000000000000";
--X40Y14, linear_LMDPL
constant Tile_X40Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X41Y14, linear_LMDPL
constant Tile_X41Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000000000000000000001010101000000000010101011010101010101010000000000000000000000000101010100000000010101010000100010001000100000000101010101111111111111111000000000000000000000000000000001111111111111111";
--X42Y14, nonlinear_LMDPL
constant Tile_X42Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000101010100000000000000000000000000000000000000000000000001001100110011001";
--X43Y14, linear_LMDPL
constant Tile_X43Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000011001100110011000000000000000001100110011001100";
--X44Y14, linear_LMDPL
constant Tile_X44Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001000100010001000";
--X45Y14, nonlinear_LMDPL
constant Tile_X45Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000001010101010101010000000000000000000000000101010100000000000000000010101010101010100000000101010100110011001100110000000000000000010101010101010100000000000000000";
--X46Y14, linear_LMDPL
constant Tile_X46Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X47Y14, linear_LMDPL
constant Tile_X47Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X48Y14, nonlinear_LMDPL
constant Tile_X48Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110101010100000000000100010001000100000000101010100110011001100110000000000000000000000000000000000100010001000100";
--X49Y14, linear_LMDPL
constant Tile_X49Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101011111111010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X50Y14, linear_LMDPL
constant Tile_X50Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010111111110000000010101010000000000000000000000000101010101010101001010101000000000101010100000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X51Y14, nonlinear_LMDPL
constant Tile_X51Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000111111110101010100000000000000001010101000000000101010101010101000000000010001000100010000000000000000000000000000000000000000000000000000010001000100010000000000000000";
--X52Y14, linear_LMDPL
constant Tile_X52Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101010101010111111111010101000000000111111110000000000000000000000000000000001010101010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X53Y14, linear_LMDPL
constant Tile_X53Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000010101010101010100000000000000000000000000000000000000000101010100101010101010101000000000000000000000000111111111010101011111111000000001010101000000000111111110000000000000000101010100101010100000000000000000000000000000000101010100000000000000000110111011101110100000000000000001110111011101110";
--X54Y14, nonlinear_LMDPL
constant Tile_X54Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000010101010101010100000000101010101100110011001100000000000000000010001000100010000000000000000000";
--X55Y14, linear_LMDPL
constant Tile_X55Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X56Y14, linear_LMDPL
constant Tile_X56Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X57Y14, nonlinear_LMDPL
constant Tile_X57Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010101010100000000000000000001000100010001";
--X58Y14, linear_LMDPL
constant Tile_X58Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X59Y14, linear_LMDPL
constant Tile_X59Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000000000000101010111111111000000000000000000000000101010100000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000011001100110011";
--X60Y14, nonlinear_LMDPL
constant Tile_X60Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101010001000100010000000000101010100000000000000000000000000000000010001000100010000000000000000000";
--X61Y14, linear_LMDPL
constant Tile_X61Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101111111111111111000000000000000011001100110011000000000000000000";
--X62Y14, linear_LMDPL
constant Tile_X62Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010";
--X63Y14, nonlinear_LMDPL
constant Tile_X63Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X64Y14, linear_LMDPL
constant Tile_X64Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001100110011001100";
--X65Y14, linear_LMDPL
constant Tile_X65Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X66Y14, nonlinear_LMDPL
constant Tile_X66Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000010101010010101010000000010101010000000000000000001010101000000000000000000000000000000000101010101010101000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y14, linear_LMDPL
constant Tile_X67Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000101010100000000000100010001000100000000000000001100110011001100000000000000000000000000000000000011001100110011";
--X68Y14, linear_LMDPL
constant Tile_X68Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000010101010000000000101010100000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000001001100110011001000000000000000011011101110111010000000000000000";
--X69Y14, nonlinear_LMDPL
constant Tile_X69Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y14, linear_LMDPL
constant Tile_X70Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000101010100000000010101010101010100000000000000001111111111111111000000000000000000100010001000100000000000000000";
--X71Y14, linear_LMDPL
constant Tile_X71Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000001010101011111111000000000101010100000000000000000000000000000000000100010001000100000000010101010101010101010101000000000000000000000000000000000010001000100010";
--X72Y14, nonlinear_LMDPL
constant Tile_X72Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X73Y14, linear_LMDPL
constant Tile_X73Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X74Y14, linear_LMDPL
constant Tile_X74Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001100110011001100000000000000000010111011101110110000000000000000";
--X75Y14, nonlinear_LMDPL
constant Tile_X75Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X76Y14, linear_LMDPL
constant Tile_X76Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X77Y14, linear_LMDPL
constant Tile_X77Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X78Y14, ctrl_to_sec
constant Tile_X78Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y14, combined_WDDL
constant Tile_X79Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y14, combined_WDDL
constant Tile_X80Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y14, ctrl_IO
constant Tile_X81Y14_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y15, W_IO_custom
constant Tile_X0Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000001010100000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000001101010100000000000000000000000000000000000000000000";
--X1Y15, linear_LMDPL
constant Tile_X1Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101011011101110111011000000000000000011001100110011000000000000000000";
--X2Y15, linear_LMDPL
constant Tile_X2Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X3Y15, nonlinear_LMDPL
constant Tile_X3Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010100000000000000001010101000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000100010001000100";
--X4Y15, linear_LMDPL
constant Tile_X4Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000010101010010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X5Y15, linear_LMDPL
constant Tile_X5Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000101010100000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X6Y15, nonlinear_LMDPL
constant Tile_X6Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000000100010001000100000000000000000";
--X7Y15, linear_LMDPL
constant Tile_X7Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001001100110011001";
--X8Y15, linear_LMDPL
constant Tile_X8Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X9Y15, nonlinear_LMDPL
constant Tile_X9Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010001000100010011111111000000000000000000000000010001000100010000010001000100010000000000000000";
--X10Y15, linear_LMDPL
constant Tile_X10Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X11Y15, linear_LMDPL
constant Tile_X11Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000011111111000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000111011101110111000000000000000001011101110111011";
--X12Y15, nonlinear_LMDPL
constant Tile_X12Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X13Y15, linear_LMDPL
constant Tile_X13Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X14Y15, linear_LMDPL
constant Tile_X14Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X15Y15, nonlinear_LMDPL
constant Tile_X15Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010100000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000011001100110011";
--X16Y15, linear_LMDPL
constant Tile_X16Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X17Y15, linear_LMDPL
constant Tile_X17Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X18Y15, nonlinear_LMDPL
constant Tile_X18Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X19Y15, linear_LMDPL
constant Tile_X19Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X20Y15, linear_LMDPL
constant Tile_X20Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000000000000010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X21Y15, nonlinear_LMDPL
constant Tile_X21Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X22Y15, linear_LMDPL
constant Tile_X22Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X23Y15, linear_LMDPL
constant Tile_X23Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000001110111011101110000000000000000";
--X24Y15, nonlinear_LMDPL
constant Tile_X24Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000100010001000100";
--X25Y15, linear_LMDPL
constant Tile_X25Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X26Y15, linear_LMDPL
constant Tile_X26Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X27Y15, nonlinear_LMDPL
constant Tile_X27Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000000000000000011111111000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X28Y15, linear_LMDPL
constant Tile_X28Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000110101010000000000100010001000100000000000000000000000000000000000000000000000000";
--X29Y15, linear_LMDPL
constant Tile_X29Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000010101010000000000000000000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000110011001100110";
--X30Y15, nonlinear_LMDPL
constant Tile_X30Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010101010100000000000000001010101000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101000000000010101011010101000000000000000000000000000000000000000000000000000000000000100010001000111111111000000001101110111011101000000000000000000000000000000000001000100010001";
--X31Y15, linear_LMDPL
constant Tile_X31Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000101010101010101101010100000000000000000101010101010101000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X32Y15, linear_LMDPL
constant Tile_X32Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000111111111010101000000000101010100000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001011101110111011";
--X33Y15, nonlinear_LMDPL
constant Tile_X33Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100100010001000100000000000000000000000000000000000110011001100110";
--X34Y15, linear_LMDPL
constant Tile_X34Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100000000000000000101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X35Y15, linear_LMDPL
constant Tile_X35Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010010101010101010100000000000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X36Y15, nonlinear_LMDPL
constant Tile_X36Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000011001100110011";
--X37Y15, linear_LMDPL
constant Tile_X37Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X38Y15, linear_LMDPL
constant Tile_X38Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000000010001000100010";
--X39Y15, nonlinear_LMDPL
constant Tile_X39Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000001010101000100010001000100000000000000000110011001100110000000000000000000000000000000000010001000100010";
--X40Y15, linear_LMDPL
constant Tile_X40Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X41Y15, linear_LMDPL
constant Tile_X41Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000000000000101010100000000010101010000100010001000100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X42Y15, nonlinear_LMDPL
constant Tile_X42Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000100010001000100";
--X43Y15, linear_LMDPL
constant Tile_X43Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000010101011010101001010101010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X44Y15, linear_LMDPL
constant Tile_X44Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101010101010101010111111111000000001000100010001000000000000000000000100010001000100000000000000000";
--X45Y15, nonlinear_LMDPL
constant Tile_X45Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000111111110000000000000000101010100000000000000000000000000101010100000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010100000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000111011101110111";
--X46Y15, linear_LMDPL
constant Tile_X46Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001111111100000000101010100000000000000000000000000101010110101010000000001010101000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X47Y15, linear_LMDPL
constant Tile_X47Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010101010101010100000000000000000";
--X48Y15, nonlinear_LMDPL
constant Tile_X48Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000010101010101010100000000101010100110011001100110000000000000000001000100010001000000000000000000";
--X49Y15, linear_LMDPL
constant Tile_X49Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000100010001000100000000000000001011101110111011000000000000000000000000000000000010001000100010";
--X50Y15, linear_LMDPL
constant Tile_X50Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X51Y15, nonlinear_LMDPL
constant Tile_X51Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010101010100000000010101010000000000000000000000000000000000101010111111111000000000101010100000000101010101010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X52Y15, linear_LMDPL
constant Tile_X52Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000101010110101010000000000000000000000000000000001010101001010101000000000000000000000000010001000100010000000000000000000000000000000000110111011101110110101010101010100000000000000000";
--X53Y15, linear_LMDPL
constant Tile_X53Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000111111111010101000000000101010101010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X54Y15, nonlinear_LMDPL
constant Tile_X54Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101001010101010101010101010100000000000000000110011001100110000000000000000010001000100010000000000000000000";
--X55Y15, linear_LMDPL
constant Tile_X55Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X56Y15, linear_LMDPL
constant Tile_X56Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000001010101000000000000000000000000000000000000000000101010100000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X57Y15, nonlinear_LMDPL
constant Tile_X57Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X58Y15, linear_LMDPL
constant Tile_X58Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X59Y15, linear_LMDPL
constant Tile_X59Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000011111111000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X60Y15, nonlinear_LMDPL
constant Tile_X60Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X61Y15, linear_LMDPL
constant Tile_X61Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010101011111111100000000000000000000000000000000000000000000000001010101101010100000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000010101010111011101110111000000000000000000000000000000000101010101010101";
--X62Y15, linear_LMDPL
constant Tile_X62Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010101010110101010000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X63Y15, nonlinear_LMDPL
constant Tile_X63Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010101010100000000010101011110111011101110000000000000000010101010101010100000000000000000";
--X64Y15, linear_LMDPL
constant Tile_X64Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010101111111101010101101010101111111100000000000000001010101000000000000000000000000000000000000000000000000000000000111111110101010100000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X65Y15, linear_LMDPL
constant Tile_X65Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000011111111000000000000000011111111000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000111011101110111000000000000000000000000000000000001000100010001";
--X66Y15, nonlinear_LMDPL
constant Tile_X66Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X67Y15, linear_LMDPL
constant Tile_X67Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X68Y15, linear_LMDPL
constant Tile_X68Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000111111111111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000000000000000000000000000000000000000000000000000111011101110111";
--X69Y15, nonlinear_LMDPL
constant Tile_X69Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000100010001000100000000101010100110011001100110000000000000000000000000000000000010001000100010";
--X70Y15, linear_LMDPL
constant Tile_X70Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X71Y15, linear_LMDPL
constant Tile_X71Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000010101010101010100000000000000001001100110011001000000000000000000100010001000100000000000000000";
--X72Y15, nonlinear_LMDPL
constant Tile_X72Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X73Y15, linear_LMDPL
constant Tile_X73Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000010101010101010100000000101010101000100010001000000000000000000011011101110111010000000000000000";
--X74Y15, linear_LMDPL
constant Tile_X74Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000000000000000000000000000000000000";
--X75Y15, nonlinear_LMDPL
constant Tile_X75Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X76Y15, linear_LMDPL
constant Tile_X76Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000101010101100110011001100000000000000000010101010101010100000000000000000";
--X77Y15, linear_LMDPL
constant Tile_X77Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X78Y15, ctrl_to_sec
constant Tile_X78Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y15, combined_WDDL
constant Tile_X79Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y15, combined_WDDL
constant Tile_X80Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y15, ctrl_IO
constant Tile_X81Y15_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y16, W_IO_custom
constant Tile_X0Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010100000000000000000000000000000000000000001111111110000000010111111111000000000000000000000000";
--X1Y16, linear_LMDPL
constant Tile_X1Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000010101010101010101110111011101110000000000000000";
--X2Y16, linear_LMDPL
constant Tile_X2Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000000000000000000000000000000000000";
--X3Y16, nonlinear_LMDPL
constant Tile_X3Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010101010100000000101010100001000100010001000000000000000010011001100110010000000000000000";
--X4Y16, linear_LMDPL
constant Tile_X4Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000010101010000000010101010010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X5Y16, linear_LMDPL
constant Tile_X5Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111101010101010001000100010000000000000000000000000000000000010101010101010101000100010001000000000000000000";
--X6Y16, nonlinear_LMDPL
constant Tile_X6Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X7Y16, linear_LMDPL
constant Tile_X7Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X8Y16, linear_LMDPL
constant Tile_X8Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000101010101010101011101110111011100000000000000000";
--X9Y16, nonlinear_LMDPL
constant Tile_X9Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111010101010101010100000000101010101001100110011001000000000000000011001100110011000000000000000000";
--X10Y16, linear_LMDPL
constant Tile_X10Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101011111111101010100000000000000000101010100000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X11Y16, linear_LMDPL
constant Tile_X11Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001011101110111011";
--X12Y16, nonlinear_LMDPL
constant Tile_X12Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000001010101000100010001000100000000000000001001100110011001000000000000000000000000000000000001000100010001";
--X13Y16, linear_LMDPL
constant Tile_X13Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001000100010001000";
--X14Y16, linear_LMDPL
constant Tile_X14Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010111111110000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000000000000000000";
--X15Y16, nonlinear_LMDPL
constant Tile_X15Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000010001000100010";
--X16Y16, linear_LMDPL
constant Tile_X16Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X17Y16, linear_LMDPL
constant Tile_X17Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100";
--X18Y16, nonlinear_LMDPL
constant Tile_X18Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000001111111111111111000000000000000000000000000000000011001100110011";
--X19Y16, linear_LMDPL
constant Tile_X19Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X20Y16, linear_LMDPL
constant Tile_X20Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X21Y16, nonlinear_LMDPL
constant Tile_X21Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000010101010000100010001000100000000010101011110111011101110000000000000000000000000000000000011001100110011";
--X22Y16, linear_LMDPL
constant Tile_X22Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000";
--X23Y16, linear_LMDPL
constant Tile_X23Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X24Y16, nonlinear_LMDPL
constant Tile_X24Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X25Y16, linear_LMDPL
constant Tile_X25Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X26Y16, linear_LMDPL
constant Tile_X26Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X27Y16, nonlinear_LMDPL
constant Tile_X27Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X28Y16, linear_LMDPL
constant Tile_X28Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000100010001000100";
--X29Y16, linear_LMDPL
constant Tile_X29Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000101010100000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000011001100110011";
--X30Y16, nonlinear_LMDPL
constant Tile_X30Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010100000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y16, linear_LMDPL
constant Tile_X31Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000001010101000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000101010100101010100000000101010100000000000000000101010100000000010101010000000000000000000000000010001000100010000000000000000000000000000000000010101010101010100000000000000000000000000000000";
--X32Y16, linear_LMDPL
constant Tile_X32Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101010101010101010100000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X33Y16, nonlinear_LMDPL
constant Tile_X33Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000100010001000100";
--X34Y16, linear_LMDPL
constant Tile_X34Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000101010101010101";
--X35Y16, linear_LMDPL
constant Tile_X35Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111111111110000000000000000101010100000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001010101010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X36Y16, nonlinear_LMDPL
constant Tile_X36Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101010101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y16, linear_LMDPL
constant Tile_X37Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001111111100000000000000000000000001010101010001000100010000000000000000000000000000000000100010001000100001110111011101110000000000000000";
--X38Y16, linear_LMDPL
constant Tile_X38Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000000000000010101010000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000110011001100110";
--X39Y16, nonlinear_LMDPL
constant Tile_X39Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000010101010000000001010101000100010001000100000000101010100011001100110011000000000000000000000000000000000010001000100010";
--X40Y16, linear_LMDPL
constant Tile_X40Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000101010101010101000000000000000001010101001010101000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X41Y16, linear_LMDPL
constant Tile_X41Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X42Y16, nonlinear_LMDPL
constant Tile_X42Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000001010101000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000010001000100010";
--X43Y16, linear_LMDPL
constant Tile_X43Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010111111111000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X44Y16, linear_LMDPL
constant Tile_X44Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X45Y16, nonlinear_LMDPL
constant Tile_X45Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000010101011110111011101110000000000000000000000000000000000000000000000000";
--X46Y16, linear_LMDPL
constant Tile_X46Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001010101010101010";
--X47Y16, linear_LMDPL
constant Tile_X47Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X48Y16, nonlinear_LMDPL
constant Tile_X48Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000010101010101010110011001100110010000000000000000";
--X49Y16, linear_LMDPL
constant Tile_X49Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010010101010101010100000000010101011000100010001000000000000000000000000000000000000000000000000000";
--X50Y16, linear_LMDPL
constant Tile_X50Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000101010101010101010101010000000000000000000000000010101010000000010101010010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X51Y16, nonlinear_LMDPL
constant Tile_X51Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000101010110101010101010100000000000000000000000000000000000000000010101011010101000000000000000000101010100000000000000001010101011111111010001000100010000000000000000000000000000000000011101110111011110001000100010000000000000000000";
--X52Y16, linear_LMDPL
constant Tile_X52Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X53Y16, linear_LMDPL
constant Tile_X53Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101111111100000000101010100000000000000000000000001111111100000000010101010101010100000000000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100";
--X54Y16, nonlinear_LMDPL
constant Tile_X54Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101010101001010101000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010101010101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X55Y16, linear_LMDPL
constant Tile_X55Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X56Y16, linear_LMDPL
constant Tile_X56Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000001010101001010101010101010101010100000000000000000001000100010001000000000000000000000000000000000000000000000000";
--X57Y16, nonlinear_LMDPL
constant Tile_X57Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000101010100101010101010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000101010100110011001100110000000000000000001010101010101010000000000000000";
--X58Y16, linear_LMDPL
constant Tile_X58Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X59Y16, linear_LMDPL
constant Tile_X59Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000010001000100010000000000101010100000000000000000100010001000100010101010101010100000000000000000";
--X60Y16, nonlinear_LMDPL
constant Tile_X60Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y16, linear_LMDPL
constant Tile_X61Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010101010101000100010001000100000000101010100100010001000100000000000000000000000000000000000100010001000100";
--X62Y16, linear_LMDPL
constant Tile_X62Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111110101010000000001010101000000000000000001010101011111111010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X63Y16, nonlinear_LMDPL
constant Tile_X63Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000101110111011101100000000000000000101010101010101";
--X64Y16, linear_LMDPL
constant Tile_X64Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101011010101011111111000000000000000000000000000000000000000001010101101010100000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000101010101101010101100110011001100000000000000000000000000000000001111111111111111";
--X65Y16, linear_LMDPL
constant Tile_X65Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000111011101110111";
--X66Y16, nonlinear_LMDPL
constant Tile_X66Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010001000100010000000000101010100000000000000000001100110011001101010101010101010000000000000000";
--X67Y16, linear_LMDPL
constant Tile_X67Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000010101010101010101111111100000000000000001111111110101010000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X68Y16, linear_LMDPL
constant Tile_X68Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010001010101000000000000000000000000101010101010101001110111011101110000000000000000";
--X69Y16, nonlinear_LMDPL
constant Tile_X69Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010110101010010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X70Y16, linear_LMDPL
constant Tile_X70Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X71Y16, linear_LMDPL
constant Tile_X71Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000000000000000000";
--X72Y16, nonlinear_LMDPL
constant Tile_X72Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000001000100010001010101010101010100000000000000000";
--X73Y16, linear_LMDPL
constant Tile_X73Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X74Y16, linear_LMDPL
constant Tile_X74Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000001100110011001100000000000000000000000000000000";
--X75Y16, nonlinear_LMDPL
constant Tile_X75Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X76Y16, linear_LMDPL
constant Tile_X76Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X77Y16, linear_LMDPL
constant Tile_X77Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000001100110011001100000000000000000100010001000100";
--X78Y16, ctrl_to_sec
constant Tile_X78Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y16, combined_WDDL
constant Tile_X79Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y16, combined_WDDL
constant Tile_X80Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y16, ctrl_IO
constant Tile_X81Y16_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y17, W_IO_custom
constant Tile_X0Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000001010100000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000001101010100000000000000000000110110110110000000000000";
--X1Y17, linear_LMDPL
constant Tile_X1Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X2Y17, linear_LMDPL
constant Tile_X2Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X3Y17, nonlinear_LMDPL
constant Tile_X3Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000010001000100010000000000000000";
--X4Y17, linear_LMDPL
constant Tile_X4Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000010101010000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X5Y17, linear_LMDPL
constant Tile_X5Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111111010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001010101010101010";
--X6Y17, nonlinear_LMDPL
constant Tile_X6Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X7Y17, linear_LMDPL
constant Tile_X7Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001010101010101010";
--X8Y17, linear_LMDPL
constant Tile_X8Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X9Y17, nonlinear_LMDPL
constant Tile_X9Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001001100110011001";
--X10Y17, linear_LMDPL
constant Tile_X10Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X11Y17, linear_LMDPL
constant Tile_X11Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001110111011101110";
--X12Y17, nonlinear_LMDPL
constant Tile_X12Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000000000000010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X13Y17, linear_LMDPL
constant Tile_X13Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000110011001100110";
--X14Y17, linear_LMDPL
constant Tile_X14Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000110011001100110001010101010101010000000000000000";
--X15Y17, nonlinear_LMDPL
constant Tile_X15Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X16Y17, linear_LMDPL
constant Tile_X16Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001110111011101110";
--X17Y17, linear_LMDPL
constant Tile_X17Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X18Y17, nonlinear_LMDPL
constant Tile_X18Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y17, linear_LMDPL
constant Tile_X19Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011";
--X20Y17, linear_LMDPL
constant Tile_X20Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X21Y17, nonlinear_LMDPL
constant Tile_X21Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000011001100110011";
--X22Y17, linear_LMDPL
constant Tile_X22Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X23Y17, linear_LMDPL
constant Tile_X23Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000111111111010101010010001000100010000000000000000000000000000000000000000000000000";
--X24Y17, nonlinear_LMDPL
constant Tile_X24Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X25Y17, linear_LMDPL
constant Tile_X25Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001101110111011101";
--X26Y17, linear_LMDPL
constant Tile_X26Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X27Y17, nonlinear_LMDPL
constant Tile_X27Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000011001100110011000000000000000000101010101010101";
--X28Y17, linear_LMDPL
constant Tile_X28Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000001000100010001";
--X29Y17, linear_LMDPL
constant Tile_X29Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X30Y17, nonlinear_LMDPL
constant Tile_X30Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000101010101010101";
--X31Y17, linear_LMDPL
constant Tile_X31Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101000000000111111110000000000000000000000001111111100000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X32Y17, linear_LMDPL
constant Tile_X32Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100101010100000000000000001010101010101010101010100000000000000000000000001111111100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X33Y17, nonlinear_LMDPL
constant Tile_X33Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X34Y17, linear_LMDPL
constant Tile_X34Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001110111011101110000000000000000";
--X35Y17, linear_LMDPL
constant Tile_X35Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X36Y17, nonlinear_LMDPL
constant Tile_X36Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010110101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000000100010001000100";
--X37Y17, linear_LMDPL
constant Tile_X37Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000010101010111111111010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X38Y17, linear_LMDPL
constant Tile_X38Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000000000000000000000010101010101010100000000010101010101010100000000101010101000100010001000000000000000000001010101010101010000000000000000";
--X39Y17, nonlinear_LMDPL
constant Tile_X39Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X40Y17, linear_LMDPL
constant Tile_X40Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000101010100000000000000000111111111010101000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000010101010000000000000000010001000100010000000000000000001010101010101010";
--X41Y17, linear_LMDPL
constant Tile_X41Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X42Y17, nonlinear_LMDPL
constant Tile_X42Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010010101010000000010101010101010100000000000000000101010100101010100000000000000000101010100000000000000000000000011111111000000000101010100000000010101010101010100000000101010100111011101110111000000000000000010001000100010000000000000000000";
--X43Y17, linear_LMDPL
constant Tile_X43Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X44Y17, linear_LMDPL
constant Tile_X44Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X45Y17, nonlinear_LMDPL
constant Tile_X45Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101111111100000000010101011010101000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X46Y17, linear_LMDPL
constant Tile_X46Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000001010101001010101000000000101010110101010000000000000000000000000000000000000000000000000100010001000100000000000000000000111011101110111";
--X47Y17, linear_LMDPL
constant Tile_X47Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000010101010000000000101010100000000111111110000000000000000000100010001000100000000101010100000000000000000000000000000000000000000000000001010101010101010";
--X48Y17, nonlinear_LMDPL
constant Tile_X48Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000001010101000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000101010101010101";
--X49Y17, linear_LMDPL
constant Tile_X49Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X50Y17, linear_LMDPL
constant Tile_X50Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000010101010000000001010101101010100000000000000000000000001010101000000000101010100000000001010101000000000000000000000000000000000101010110101010000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X51Y17, nonlinear_LMDPL
constant Tile_X51Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100101010100000000000000000101010100000000101010100000000001010101010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000100010001000100000000101010100110011001100110000000000000000000000000000000000000000000000000";
--X52Y17, linear_LMDPL
constant Tile_X52Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000010101010000000000000000111111110000000000000000101010101010101000000000101010100101010100000000000000000101010101010101000000000101010110101010000000000000000011111111000000000000000000000000000000000000000000000000000000000100010001000100";
--X53Y17, linear_LMDPL
constant Tile_X53Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X54Y17, nonlinear_LMDPL
constant Tile_X54Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000101010110101010000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000001000100010001000000000000000000";
--X55Y17, linear_LMDPL
constant Tile_X55Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110011011101110111010000000000000000";
--X56Y17, linear_LMDPL
constant Tile_X56Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000010011001100110010000000000000000";
--X57Y17, nonlinear_LMDPL
constant Tile_X57Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000000000000000000000";
--X58Y17, linear_LMDPL
constant Tile_X58Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101011111111100000000101010100000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000101010100000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010";
--X59Y17, linear_LMDPL
constant Tile_X59Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100000000000000000010101010000000000000000000000001111111101010101000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X60Y17, nonlinear_LMDPL
constant Tile_X60Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000101010100000000000000001010101000000000000000000101010101010101000000000000000000000000000000001111111100000000000000000101010101010101000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000011001100110011001000100010001000000000000000000";
--X61Y17, linear_LMDPL
constant Tile_X61Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000010001000100010000000000101010100000000000000000000000000000000010101010101010100000000000000000";
--X62Y17, linear_LMDPL
constant Tile_X62Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000001010101000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X63Y17, nonlinear_LMDPL
constant Tile_X63Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X64Y17, linear_LMDPL
constant Tile_X64Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000001010101000000000000000000000000101010100000000001010101101010100000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X65Y17, linear_LMDPL
constant Tile_X65Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X66Y17, nonlinear_LMDPL
constant Tile_X66Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y17, linear_LMDPL
constant Tile_X67Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000010101010101010100000000000000000000000001111111110101010101010100000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X68Y17, linear_LMDPL
constant Tile_X68Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101010001000100010000000000010101010000000000000000100010001000100010001000100010000000000000000000";
--X69Y17, nonlinear_LMDPL
constant Tile_X69Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y17, linear_LMDPL
constant Tile_X70Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000010101011100110011001100000000000000000000000000000000001010101010101010";
--X71Y17, linear_LMDPL
constant Tile_X71Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000001000100010001000000000000000001000100010001000";
--X72Y17, nonlinear_LMDPL
constant Tile_X72Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X73Y17, linear_LMDPL
constant Tile_X73Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111101010100000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010";
--X74Y17, linear_LMDPL
constant Tile_X74Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000000010001000100010";
--X75Y17, nonlinear_LMDPL
constant Tile_X75Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010101010101010100000000101010101011101110111011000000000000000000000000000000000000000000000000";
--X76Y17, linear_LMDPL
constant Tile_X76Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100010001000100010000000000000000000000000000000000101010101010101";
--X77Y17, linear_LMDPL
constant Tile_X77Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X78Y17, ctrl_to_sec
constant Tile_X78Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y17, combined_WDDL
constant Tile_X79Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y17, combined_WDDL
constant Tile_X80Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y17, ctrl_IO
constant Tile_X81Y17_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y18, W_IO_custom
constant Tile_X0Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000110110110110";
--X1Y18, linear_LMDPL
constant Tile_X1Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X2Y18, linear_LMDPL
constant Tile_X2Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000010001000100010000000000111111110000000000000000101110111011101100000000000000000000000000000000";
--X3Y18, nonlinear_LMDPL
constant Tile_X3Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000011011101110111010000000000000000";
--X4Y18, linear_LMDPL
constant Tile_X4Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000101010100000000000000000111111111010101000000000000000000000000000000000000000000101010110101010000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X5Y18, linear_LMDPL
constant Tile_X5Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X6Y18, nonlinear_LMDPL
constant Tile_X6Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010011001100110010000000000000000";
--X7Y18, linear_LMDPL
constant Tile_X7Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X8Y18, linear_LMDPL
constant Tile_X8Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010101010000000011111111010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X9Y18, nonlinear_LMDPL
constant Tile_X9Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000101010101111111111111111000000000000000010101010101010100000000000000000";
--X10Y18, linear_LMDPL
constant Tile_X10Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000110011001100110000000000000000";
--X11Y18, linear_LMDPL
constant Tile_X11Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000101010101010101011111111010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X12Y18, nonlinear_LMDPL
constant Tile_X12Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000001010101010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X13Y18, linear_LMDPL
constant Tile_X13Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X14Y18, linear_LMDPL
constant Tile_X14Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X15Y18, nonlinear_LMDPL
constant Tile_X15Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000001011101110111011";
--X16Y18, linear_LMDPL
constant Tile_X16Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X17Y18, linear_LMDPL
constant Tile_X17Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X18Y18, nonlinear_LMDPL
constant Tile_X18Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000001101110111011101000000000000000000010001000100010000000000000000";
--X19Y18, linear_LMDPL
constant Tile_X19Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X20Y18, linear_LMDPL
constant Tile_X20Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000011111111010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X21Y18, nonlinear_LMDPL
constant Tile_X21Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000011001100110011";
--X22Y18, linear_LMDPL
constant Tile_X22Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110000000010101010010101010101010100000000101010100000000000000000000000000000000001110111011101110000000000000000";
--X23Y18, linear_LMDPL
constant Tile_X23Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000111111110100010001000100000000000000000011011101110111010000000000000000";
--X24Y18, nonlinear_LMDPL
constant Tile_X24Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X25Y18, linear_LMDPL
constant Tile_X25Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001010101010101010000000000000000010011001100110010000000000000000";
--X26Y18, linear_LMDPL
constant Tile_X26Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X27Y18, nonlinear_LMDPL
constant Tile_X27Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101011010101010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100110011001100100000000000000000010001000100010";
--X28Y18, linear_LMDPL
constant Tile_X28Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000001111111111111111000000000000000011101110111011100000000000000000";
--X29Y18, linear_LMDPL
constant Tile_X29Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X30Y18, nonlinear_LMDPL
constant Tile_X30Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101010101011111111100000000000000000000000000000000000000000000000001010101010101010000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000011111111000100010001000100000000000000001111111111111111000000000000000000000000000000000010001000100010";
--X31Y18, linear_LMDPL
constant Tile_X31Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000111111111010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X32Y18, linear_LMDPL
constant Tile_X32Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101010101010101010100101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001111111111111111";
--X33Y18, nonlinear_LMDPL
constant Tile_X33Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000000010001000100010";
--X34Y18, linear_LMDPL
constant Tile_X34Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X35Y18, linear_LMDPL
constant Tile_X35Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X36Y18, nonlinear_LMDPL
constant Tile_X36Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000001010101111111110000000000000000000000000101010100000000000000000000000000000000000100010001000100000000101010101000100010001000000000000000000000000000000000000010001000100010";
--X37Y18, linear_LMDPL
constant Tile_X37Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000001111111100000000101010101111111100000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X38Y18, linear_LMDPL
constant Tile_X38Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000010101010010101011010101000000000010001000100010000000000000000000000000000000000110111011101110101110111011101110000000000000000";
--X39Y18, nonlinear_LMDPL
constant Tile_X39Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X40Y18, linear_LMDPL
constant Tile_X40Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101000000000111111110000000000000000000000000000000010101010101010100000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X41Y18, linear_LMDPL
constant Tile_X41Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000111111110000000010101010010001000100010000000000101010100000000000000000101010101010101011001100110011000000000000000000";
--X42Y18, nonlinear_LMDPL
constant Tile_X42Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100101010110101010010101010000000000000000000000000000000001010101000000001010101000000000000000000000000011111111000000000000000001010101000100010001000100000000101010100001000100010001000000000000000000000000000000001100110011001100";
--X43Y18, linear_LMDPL
constant Tile_X43Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010111111111000000000000000010101010000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000101010101010101";
--X44Y18, linear_LMDPL
constant Tile_X44Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101000000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000001111111111111111000000000000000000000000000000001111111111111111";
--X45Y18, nonlinear_LMDPL
constant Tile_X45Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000010001000100010";
--X46Y18, linear_LMDPL
constant Tile_X46Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000101010100000000001010101000000000000000001010101000000000000000000000000000000000000000010101010000100010001000100000000111111111000100010001000000000000000000000000000000000000000000000000000";
--X47Y18, linear_LMDPL
constant Tile_X47Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110101010110101010000000000000000000000000000000000000000001010101010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X48Y18, nonlinear_LMDPL
constant Tile_X48Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000101110111011101110001000100010000000000000000000";
--X49Y18, linear_LMDPL
constant Tile_X49Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000101010100101010100000000101010100000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000001001100110011001";
--X50Y18, linear_LMDPL
constant Tile_X50Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010101010100000000010101010000000000000000000000000000000001010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X51Y18, nonlinear_LMDPL
constant Tile_X51Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X52Y18, linear_LMDPL
constant Tile_X52Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000101010100000000001010101000000000000000000000000000000001010101010101010101010101010101000000000000000000000000011111111000000000101010110101010000100010001000100000000000000000101010101010101000000000000000000000000000000000000000000000000";
--X53Y18, linear_LMDPL
constant Tile_X53Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000010101010000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000101010100000000010001000100010000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X54Y18, nonlinear_LMDPL
constant Tile_X54Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000000000000000000000";
--X55Y18, linear_LMDPL
constant Tile_X55Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000101010100000000000000000000000000000000111111110000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X56Y18, linear_LMDPL
constant Tile_X56Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X57Y18, nonlinear_LMDPL
constant Tile_X57Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010110101010000000000000000000000000010101011010101000000000010101011010101000000000000000000000000000000000000000001010101000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X58Y18, linear_LMDPL
constant Tile_X58Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010101010101010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X59Y18, linear_LMDPL
constant Tile_X59Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000010101010101010100000000111111110000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000101010100000000010101010101010100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X60Y18, nonlinear_LMDPL
constant Tile_X60Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y18, linear_LMDPL
constant Tile_X61Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000010101010000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010111111111000100010001000100000000101010100100010001000100000000000000000000000000000000001000100010001000";
--X62Y18, linear_LMDPL
constant Tile_X62Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000000000001111111100000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X63Y18, nonlinear_LMDPL
constant Tile_X63Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000010001000100010";
--X64Y18, linear_LMDPL
constant Tile_X64Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000000000000101010100000000010101010000000001010101000000000101010100000000011111111000000000000000001010101000000000101010100000000000000000000000000000000101010100000000000000000100110011001100100000000000000000010001000100010";
--X65Y18, linear_LMDPL
constant Tile_X65Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010111111111000000000000000000000000000000000000000000000000110111011101110100000000000000000010001000100010";
--X66Y18, nonlinear_LMDPL
constant Tile_X66Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000001100110011001100100010001000100000000000000000";
--X67Y18, linear_LMDPL
constant Tile_X67Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000101010110101010101010100000000000000000000000000000000010101010111111110000000010101010000000000000000011111111000000001010101001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101";
--X68Y18, linear_LMDPL
constant Tile_X68Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010101010101000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X69Y18, nonlinear_LMDPL
constant Tile_X69Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000010101010010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X70Y18, linear_LMDPL
constant Tile_X70Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011010001000100010000000000000000000";
--X71Y18, linear_LMDPL
constant Tile_X71Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000010001000100010000000000101010100000000000000000010001000100010010001000100010000000000000000000";
--X72Y18, nonlinear_LMDPL
constant Tile_X72Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X73Y18, linear_LMDPL
constant Tile_X73Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000000101010101010101";
--X74Y18, linear_LMDPL
constant Tile_X74Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001000100010001000";
--X75Y18, nonlinear_LMDPL
constant Tile_X75Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000110011001100110000010001000100010000000000000000";
--X76Y18, linear_LMDPL
constant Tile_X76Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X77Y18, linear_LMDPL
constant Tile_X77Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000100010001000100000000101010101001100110011001000000000000000000000000000000000100010001000100";
--X78Y18, ctrl_to_sec
constant Tile_X78Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y18, combined_WDDL
constant Tile_X79Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y18, combined_WDDL
constant Tile_X80Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y18, ctrl_IO
constant Tile_X81Y18_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y19, W_IO_custom
constant Tile_X0Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000001010100000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000";
--X1Y19, linear_LMDPL
constant Tile_X1Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011111111100000000000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X2Y19, linear_LMDPL
constant Tile_X2Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001011101110111011";
--X3Y19, nonlinear_LMDPL
constant Tile_X3Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X4Y19, linear_LMDPL
constant Tile_X4Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010101010101010101010010101010101010100000000000000001001100110011001000000000000000000100010001000100000000000000000";
--X5Y19, linear_LMDPL
constant Tile_X5Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001001100110011001";
--X6Y19, nonlinear_LMDPL
constant Tile_X6Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001001100110011001000000000000000000100010001000100000000000000000";
--X7Y19, linear_LMDPL
constant Tile_X7Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X8Y19, linear_LMDPL
constant Tile_X8Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000101010100000000010101010000000001010101000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000101010101010101";
--X9Y19, nonlinear_LMDPL
constant Tile_X9Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000011001100110011";
--X10Y19, linear_LMDPL
constant Tile_X10Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000011111111111111110000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001111111111111111";
--X11Y19, linear_LMDPL
constant Tile_X11Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X12Y19, nonlinear_LMDPL
constant Tile_X12Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X13Y19, linear_LMDPL
constant Tile_X13Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111111111110000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X14Y19, linear_LMDPL
constant Tile_X14Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010111111110000000000000000000000000000000000000000000000001010101011111111010001000100010000000000010101010000000000000000101010101010101000100010001000100000000000000000";
--X15Y19, nonlinear_LMDPL
constant Tile_X15Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000100100010001000100000000000000000";
--X16Y19, linear_LMDPL
constant Tile_X16Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010110101010000000000000000000000000000000000000000000000000111111111010101000000000000000001010101000000000010101011010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X17Y19, linear_LMDPL
constant Tile_X17Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000101010101010101000000000000000000100010001000100000000000000000";
--X18Y19, nonlinear_LMDPL
constant Tile_X18Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X19Y19, linear_LMDPL
constant Tile_X19Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X20Y19, linear_LMDPL
constant Tile_X20Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000001010101010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X21Y19, nonlinear_LMDPL
constant Tile_X21Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000100010001000100";
--X22Y19, linear_LMDPL
constant Tile_X22Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X23Y19, linear_LMDPL
constant Tile_X23Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000010101010000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X24Y19, nonlinear_LMDPL
constant Tile_X24Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000101010101010101";
--X25Y19, linear_LMDPL
constant Tile_X25Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001101110111011101000000000000000000000000000000001100110011001100";
--X26Y19, linear_LMDPL
constant Tile_X26Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X27Y19, nonlinear_LMDPL
constant Tile_X27Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X28Y19, linear_LMDPL
constant Tile_X28Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000100010001000100";
--X29Y19, linear_LMDPL
constant Tile_X29Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X30Y19, nonlinear_LMDPL
constant Tile_X30Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y19, linear_LMDPL
constant Tile_X31Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000101010101010101";
--X32Y19, linear_LMDPL
constant Tile_X32Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000001010101010101010101010100000000000000000000000000000000000000000111111110000000000000000000100010001000100000000111111110000000000000000000000000000000000000000000000000000000000000000";
--X33Y19, nonlinear_LMDPL
constant Tile_X33Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001110111011101110000000000000000001000100010001000000000000000000";
--X34Y19, linear_LMDPL
constant Tile_X34Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000101010100000000000000000000000001010101010101010010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000111011101110111";
--X35Y19, linear_LMDPL
constant Tile_X35Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000011001100110011000000000000000000";
--X36Y19, nonlinear_LMDPL
constant Tile_X36Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000000000000000000";
--X37Y19, linear_LMDPL
constant Tile_X37Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000101010110101010101010101010101000000000000000000000000000000000111111110000000001010101010001000100010000000000000000000000000000000000010001000100010001010101010101010000000000000000";
--X38Y19, linear_LMDPL
constant Tile_X38Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000111111110000000000000000000100010001000100000000101010100100010001000100000000000000000000000000000000001000100010001000";
--X39Y19, nonlinear_LMDPL
constant Tile_X39Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101110111011101110001000100010000000000000000000";
--X40Y19, linear_LMDPL
constant Tile_X40Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000101010100000000000000000001000100010001000000000000000001010101010101010";
--X41Y19, linear_LMDPL
constant Tile_X41Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010010001000100010000000000010101010000000000000000001000100010001011001100110011000000000000000000";
--X42Y19, nonlinear_LMDPL
constant Tile_X42Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000101010100000000000000001010101001010101000000001010101010101010010101010000000000000000101010100000000000000000010101010000000000000000000000000000000000000000010101010000000011111111010001000100010000000000101010100000000000000000001000100010001010011001100110010000000000000000";
--X43Y19, linear_LMDPL
constant Tile_X43Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000011111111000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000110011001100110000000000000000000100010001000100";
--X44Y19, linear_LMDPL
constant Tile_X44Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000000000000010101010101010100000000000000000000000010101010000000000000000011111111101010100000000010101010010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X45Y19, nonlinear_LMDPL
constant Tile_X45Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010101010100000000000000000010101011010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X46Y19, linear_LMDPL
constant Tile_X46Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000010101010000000000101010110101010000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000111011101110111";
--X47Y19, linear_LMDPL
constant Tile_X47Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000001010101010101010000000000000000010101010000000000000000000000000101010100101010110101010000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000111011101110111";
--X48Y19, nonlinear_LMDPL
constant Tile_X48Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001001100110011001";
--X49Y19, linear_LMDPL
constant Tile_X49Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000100010001000100000000010101011000100010001000000000000000000000000000000000000000000000000000";
--X50Y19, linear_LMDPL
constant Tile_X50Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000001010101010101010101010100000000000000000000000000000000000000000111111110101010110101010000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X51Y19, nonlinear_LMDPL
constant Tile_X51Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010001000100010000000000101010100000000000000000011101110111011101110111011101110000000000000000";
--X52Y19, linear_LMDPL
constant Tile_X52Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000011111111000000001010101000000000101010100000000001010101000000000000000000000000101010101010101010101010101010101010101000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X53Y19, linear_LMDPL
constant Tile_X53Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101010101010111111110000000010101010000000000000000000000000010101010101010100000000010101010101010100000000000000000111011101110111000000000000000001000100010001000000000000000000";
--X54Y19, nonlinear_LMDPL
constant Tile_X54Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001100110011001100";
--X55Y19, linear_LMDPL
constant Tile_X55Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000101010110101010111111110000000000000000000000001010101010101010111111111010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001111111111111111";
--X56Y19, linear_LMDPL
constant Tile_X56Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000101010100000000000000001010101000000000010101010000000000000000000000000000000000000000010101011010101000000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X57Y19, nonlinear_LMDPL
constant Tile_X57Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000010101011111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000101010101010101000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100110011001100110000000000000000000000000000000000000000000000000";
--X58Y19, linear_LMDPL
constant Tile_X58Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101001010101101010100000000000000000000000000000000010101010101010100000000000000000010101010101010100000000101010101010101010101010000000000000000000000000000000000000000000000000";
--X59Y19, linear_LMDPL
constant Tile_X59Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101010101011010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000111011101110111";
--X60Y19, nonlinear_LMDPL
constant Tile_X60Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101011010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X61Y19, linear_LMDPL
constant Tile_X61Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000101010100000000101010100000000000000000000000000101010100000000010101010000000000000000000000001010101010101010000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010100000000000000000011101110111011100000000000000000100010001000100";
--X62Y19, linear_LMDPL
constant Tile_X62Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X63Y19, nonlinear_LMDPL
constant Tile_X63Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010001000100010000000000101010100000000000000000011001100110011000100010001000100000000000000000";
--X64Y19, linear_LMDPL
constant Tile_X64Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010101010101000000000000000001010101000000000101010100000000010101010101010101010101000000000000000001010101000000000010101010101010100000000010101010010001000100010000000000000000000000000000000000000000000000000";
--X65Y19, linear_LMDPL
constant Tile_X65Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000010101010000000001111111100000000000000000000000000000000101010101010101000000000000000000000000011111111000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000110011001100110000000000000000001111111111111111";
--X66Y19, nonlinear_LMDPL
constant Tile_X66Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y19, linear_LMDPL
constant Tile_X67Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101001010101101010100000000000000000000000000000000010101010111111110000000010101010000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X68Y19, linear_LMDPL
constant Tile_X68Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101010101010";
--X69Y19, nonlinear_LMDPL
constant Tile_X69Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y19, linear_LMDPL
constant Tile_X70Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000000100010001000110001000100010000000000000000000";
--X71Y19, linear_LMDPL
constant Tile_X71Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010010101010000000000000000000000000000000011111111101010100000000000000000001000100010001000000000000000000100010001000100";
--X72Y19, nonlinear_LMDPL
constant Tile_X72Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101011010101000000000010001000100010000000000000000000000000000000000100110011001100101000100010001000000000000000000";
--X73Y19, linear_LMDPL
constant Tile_X73Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000101010100000000000000000110011001100110010011001100110010000000000000000";
--X74Y19, linear_LMDPL
constant Tile_X74Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011";
--X75Y19, nonlinear_LMDPL
constant Tile_X75Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101111111100000000010001000100010000000000101010100000000000000000100010001000100000110011001100110000000000000000";
--X76Y19, linear_LMDPL
constant Tile_X76Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000010001000100010000000000000000001001100110011001";
--X77Y19, linear_LMDPL
constant Tile_X77Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X78Y19, ctrl_to_sec
constant Tile_X78Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y19, combined_WDDL
constant Tile_X79Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X80Y19, combined_WDDL
constant Tile_X80Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000001010000000000000000000000000000000000000000000000000";
--X81Y19, ctrl_IO
constant Tile_X81Y19_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y20, W_IO_custom
constant Tile_X0Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000";
--X1Y20, linear_LMDPL
constant Tile_X1Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X2Y20, linear_LMDPL
constant Tile_X2Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X3Y20, nonlinear_LMDPL
constant Tile_X3Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000010001000100010000010001000100010000000000000000";
--X4Y20, linear_LMDPL
constant Tile_X4Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000000000000000000001100110011001100000000000000000";
--X5Y20, linear_LMDPL
constant Tile_X5Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000001111111101010101010001000100010000000000010101010000000000000000101010101010101010111011101110110000000000000000";
--X6Y20, nonlinear_LMDPL
constant Tile_X6Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001101110111011101000000000000000011001100110011000000000000000000";
--X7Y20, linear_LMDPL
constant Tile_X7Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110111011101110101000100010001000000000000000000";
--X8Y20, linear_LMDPL
constant Tile_X8Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000001010101010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X9Y20, nonlinear_LMDPL
constant Tile_X9Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010001000100010000000000000000001011101110111011";
--X10Y20, linear_LMDPL
constant Tile_X10Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100000000011111111000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X11Y20, linear_LMDPL
constant Tile_X11Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010101010000000010101010101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X12Y20, nonlinear_LMDPL
constant Tile_X12Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X13Y20, linear_LMDPL
constant Tile_X13Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101011111111100000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X14Y20, linear_LMDPL
constant Tile_X14Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000001010101010101010101010100000000000000000000000001010101010101010010101010000000000000000000000000000000000000000010101011010101000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X15Y20, nonlinear_LMDPL
constant Tile_X15Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000001111111100000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X16Y20, linear_LMDPL
constant Tile_X16Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000001010101000000000101010101010101001010101000000000000000000000000000000001010101001010101010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X17Y20, linear_LMDPL
constant Tile_X17Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000101010100000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X18Y20, nonlinear_LMDPL
constant Tile_X18Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000011111111000000000000000000000000010101010000000010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X19Y20, linear_LMDPL
constant Tile_X19Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000011111111000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X20Y20, linear_LMDPL
constant Tile_X20Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X21Y20, nonlinear_LMDPL
constant Tile_X21Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000001010101010101010";
--X22Y20, linear_LMDPL
constant Tile_X22Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000010101010101010100000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X23Y20, linear_LMDPL
constant Tile_X23Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000110101010101010100100010001000100000000000000000000000000000000000101010101010101";
--X24Y20, nonlinear_LMDPL
constant Tile_X24Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000101010101010101";
--X25Y20, linear_LMDPL
constant Tile_X25Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001101110111011101";
--X26Y20, linear_LMDPL
constant Tile_X26Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X27Y20, nonlinear_LMDPL
constant Tile_X27Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X28Y20, linear_LMDPL
constant Tile_X28Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X29Y20, linear_LMDPL
constant Tile_X29Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000111011101110111";
--X30Y20, nonlinear_LMDPL
constant Tile_X30Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y20, linear_LMDPL
constant Tile_X31Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000011001100110011";
--X32Y20, linear_LMDPL
constant Tile_X32Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101011111111101010100000000000000000010101010000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111011001100110011000000000000000000";
--X33Y20, nonlinear_LMDPL
constant Tile_X33Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000101010101010101";
--X34Y20, linear_LMDPL
constant Tile_X34Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X35Y20, linear_LMDPL
constant Tile_X35Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000101010100101010100000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000100010001000100001010101010101010000000000000000";
--X36Y20, nonlinear_LMDPL
constant Tile_X36Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y20, linear_LMDPL
constant Tile_X37Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000000000000101010100000000000000001010101001010101101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000100010001000100";
--X38Y20, linear_LMDPL
constant Tile_X38Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000111111110000000000000000111111110000000000000000000000000101010100000000000000000000000010101010101010100000000001010101010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X39Y20, nonlinear_LMDPL
constant Tile_X39Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010000000001010101000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000101010101010101000010001000100010000000000000000";
--X40Y20, linear_LMDPL
constant Tile_X40Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000111111110000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000000100010001000100000000000000000011011101110111010000000000000000";
--X41Y20, linear_LMDPL
constant Tile_X41Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000010101010000100010001000100000000101010100001000100010001000000000000000000000000000000001000100010001000";
--X42Y20, nonlinear_LMDPL
constant Tile_X42Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000010101010101010100000000000000000000000010101010000000000000000001010101010101010000000000000000000000000101010100000000101010100000000011111111000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000011011101110111010000000000000000";
--X43Y20, linear_LMDPL
constant Tile_X43Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111101010100000000000000000000000000000000001010101000000000000000001010101101010100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010010101011010101000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000111011101110111";
--X44Y20, linear_LMDPL
constant Tile_X44Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000011111111010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X45Y20, nonlinear_LMDPL
constant Tile_X45Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000111111110101010100000000000000000000000000000000101010100000000001010101010001000100010000000000101010100000000000000000001000100010001000010001000100010000000000000000";
--X46Y20, linear_LMDPL
constant Tile_X46Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000011111111000000000000000000000000000000000101010110101010010001000100010000000000101010100000000000000000101010101010101010001000100010000000000000000000";
--X47Y20, linear_LMDPL
constant Tile_X47Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000011111111010001000100010000000000010101010000000000000000001000100010001001000100010001000000000000000000";
--X48Y20, nonlinear_LMDPL
constant Tile_X48Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000001010101101010100000000000000000000000000000000001010101000000000101010111111111000000000000000000000000010101011010101000000000010101010101010100000000101010100001000100010001000000000000000010001000100010000000000000000000";
--X49Y20, linear_LMDPL
constant Tile_X49Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X50Y20, linear_LMDPL
constant Tile_X50Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000000000000000000000101010100000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000010001000100010";
--X51Y20, nonlinear_LMDPL
constant Tile_X51Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101011010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000100010001000100";
--X52Y20, linear_LMDPL
constant Tile_X52Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010000000000000000011111111101010100000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000001010101010101010101010100000000000000000000000000000000011111111000000000101010100000000010001000100010010101010000000000000000000000000001000100010001011001100110011000000000000000000";
--X53Y20, linear_LMDPL
constant Tile_X53Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101011111111101010101000000000000000000000000010101011010101001010101000000000000000010101010000000000000000000000000101010101010101011111111000100010001000100000000101010100010001000100010000000000000000000000000000000001010101010101010";
--X54Y20, nonlinear_LMDPL
constant Tile_X54Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000101010110101010000000000101010100000000000000000000000000000000010101010101010100000000101010100110011001100110000000000000000000100010001000100000000000000000";
--X55Y20, linear_LMDPL
constant Tile_X55Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000101010101010101010101010000000000000000000000001010101010101010010101010000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X56Y20, linear_LMDPL
constant Tile_X56Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000110011001100110011001100110011000000000000000000";
--X57Y20, nonlinear_LMDPL
constant Tile_X57Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001111111100000000010101010000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000101010100000000000100010001000100000000101010101110111011101110000000000000000000000000000000000010001000100010";
--X58Y20, linear_LMDPL
constant Tile_X58Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000010101011010101000000000010001000100010000000000000000000000000000000000100110011001100110001000100010000000000000000000";
--X59Y20, linear_LMDPL
constant Tile_X59Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000101010100000000000100010001000100000000101010100100010001000100000000000000000000000000000000000011001100110011";
--X60Y20, nonlinear_LMDPL
constant Tile_X60Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010101010101001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y20, linear_LMDPL
constant Tile_X61Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000001010101101010100000000000000000101010100000000000000000000000001010101010101010101010100101010111111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X62Y20, linear_LMDPL
constant Tile_X62Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101011010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000101010101010101";
--X63Y20, nonlinear_LMDPL
constant Tile_X63Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000010001000100010";
--X64Y20, linear_LMDPL
constant Tile_X64Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001010101000000000101010100000000010101010111111110000000010101010000000001010101000000000010001000100010000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X65Y20, linear_LMDPL
constant Tile_X65Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001101110111011101";
--X66Y20, nonlinear_LMDPL
constant Tile_X66Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y20, linear_LMDPL
constant Tile_X67Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111111111111110101010000000000000000010101010000000000000000010101010000000001010101010101010000100010001000100000000000000001101110111011101000000000000000000000000000000001100110011001100";
--X68Y20, linear_LMDPL
constant Tile_X68Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X69Y20, nonlinear_LMDPL
constant Tile_X69Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000000000000010101010000000000000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000001001100110011001";
--X70Y20, linear_LMDPL
constant Tile_X70Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101111111100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000101010101010101";
--X71Y20, linear_LMDPL
constant Tile_X71Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000010101011111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000101010100000000000000000101010101010101000000000000000000010001000100010";
--X72Y20, nonlinear_LMDPL
constant Tile_X72Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000101010100000000000000000000000000000000010001000100010000000000000000000";
--X73Y20, linear_LMDPL
constant Tile_X73Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000010101010000000000000000000000000010101010000000000000000010001000100010000000000000000000101010101010101";
--X74Y20, linear_LMDPL
constant Tile_X74Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X75Y20, nonlinear_LMDPL
constant Tile_X75Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010101010100000000101010100011001100110011000000000000000010111011101110110000000000000000";
--X76Y20, linear_LMDPL
constant Tile_X76Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010101111111110101010000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X77Y20, linear_LMDPL
constant Tile_X77Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X78Y20, ctrl_to_sec
constant Tile_X78Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y20, combined_WDDL
constant Tile_X79Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000001111000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000001000101011010000000000000000000000000100010000111011100000000";
--X80Y20, combined_WDDL
constant Tile_X80Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000101000000000000000000001000100001010111100000000000000000000101010101110111000000000";
--X81Y20, ctrl_IO
constant Tile_X81Y20_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y21, W_IO_custom
constant Tile_X0Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000001010101000000000001010100000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y21, linear_LMDPL
constant Tile_X1Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101011111111000000000000000000000000000000000000000001010101000100010001000100000000000000000000000000000000000000000000000000000000000000000101010101010101";
--X2Y21, linear_LMDPL
constant Tile_X2Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X3Y21, nonlinear_LMDPL
constant Tile_X3Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011000100010001000100000000000000000";
--X4Y21, linear_LMDPL
constant Tile_X4Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X5Y21, linear_LMDPL
constant Tile_X5Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X6Y21, nonlinear_LMDPL
constant Tile_X6Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000010001000100010";
--X7Y21, linear_LMDPL
constant Tile_X7Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X8Y21, linear_LMDPL
constant Tile_X8Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000001010101001010101000000000000000000000000000000001010101000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X9Y21, nonlinear_LMDPL
constant Tile_X9Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000010001000100010000000000000000000";
--X10Y21, linear_LMDPL
constant Tile_X10Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000111111110000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X11Y21, linear_LMDPL
constant Tile_X11Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101010101010010101010000000000000000000000001111111100000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X12Y21, nonlinear_LMDPL
constant Tile_X12Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101010101010010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X13Y21, linear_LMDPL
constant Tile_X13Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000111111110000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010111011101110110000000000000000";
--X14Y21, linear_LMDPL
constant Tile_X14Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101011010101000000000010101010101010100000000101010101100110011001100000000000000000001110111011101110000000000000000";
--X15Y21, nonlinear_LMDPL
constant Tile_X15Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110111011101110100000000000000001010101010101010";
--X16Y21, linear_LMDPL
constant Tile_X16Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000101010101010101010101010000000001111111100000000000000001010101010101010010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X17Y21, linear_LMDPL
constant Tile_X17Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101010101010010101010000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X18Y21, nonlinear_LMDPL
constant Tile_X18Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X19Y21, linear_LMDPL
constant Tile_X19Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X20Y21, linear_LMDPL
constant Tile_X20Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000101010100000000000000001010101000000000000000000000000000000000101010100000000001010101010101010101010100000000000000000100010001000100000000000000000010011001100110010000000000000000";
--X21Y21, nonlinear_LMDPL
constant Tile_X21Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000100010001000100";
--X22Y21, linear_LMDPL
constant Tile_X22Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X23Y21, linear_LMDPL
constant Tile_X23Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X24Y21, nonlinear_LMDPL
constant Tile_X24Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000010101010101010100000000010101011100110011001100000000000000000000010001000100010000000000000000";
--X25Y21, linear_LMDPL
constant Tile_X25Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X26Y21, linear_LMDPL
constant Tile_X26Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X27Y21, nonlinear_LMDPL
constant Tile_X27Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X28Y21, linear_LMDPL
constant Tile_X28Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X29Y21, linear_LMDPL
constant Tile_X29Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X30Y21, nonlinear_LMDPL
constant Tile_X30Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X31Y21, linear_LMDPL
constant Tile_X31Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X32Y21, linear_LMDPL
constant Tile_X32Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100101010100000000111111110000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000011101110111011100000000000000000";
--X33Y21, nonlinear_LMDPL
constant Tile_X33Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000000000001010101011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X34Y21, linear_LMDPL
constant Tile_X34Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000010001000100010000000000000000001110111011101110000000000000000";
--X35Y21, linear_LMDPL
constant Tile_X35Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000001111111101010101101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000001101110111011101";
--X36Y21, nonlinear_LMDPL
constant Tile_X36Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100110011001100110000000000000000010001000100010000000000000000000";
--X37Y21, linear_LMDPL
constant Tile_X37Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010110101010000000000000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X38Y21, linear_LMDPL
constant Tile_X38Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010100000000000000000000100010001000100000000101010100000000000000000000000000000000000000000000000001000100010001000";
--X39Y21, nonlinear_LMDPL
constant Tile_X39Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X40Y21, linear_LMDPL
constant Tile_X40Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X41Y21, linear_LMDPL
constant Tile_X41Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000101010100000000010101010000000000000000001010101000000000000000001010101010101010101010100000000101010100000000000000000000000000000000011001100110011000000000000000000";
--X42Y21, nonlinear_LMDPL
constant Tile_X42Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000001000100010001";
--X43Y21, linear_LMDPL
constant Tile_X43Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X44Y21, linear_LMDPL
constant Tile_X44Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001111111111111111";
--X45Y21, nonlinear_LMDPL
constant Tile_X45Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000010101011010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100101010111111111010101010101010100000000000000000001000100010001000000000000000010101010101010100000000000000000";
--X46Y21, linear_LMDPL
constant Tile_X46Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111110101010000000000000000011111111000000001010101010101010010001000100010000000000000000000000000000000000001000100010001011011101110111010000000000000000";
--X47Y21, linear_LMDPL
constant Tile_X47Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110111011101110110101010101010100000000000000000";
--X48Y21, nonlinear_LMDPL
constant Tile_X48Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000000000000101010100000000000000000000000000000000011111111101010100000000000000000101010100000000000000000000000000101010100000000000000000101010100000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000100110011001100110001000100010000000000000000000";
--X49Y21, linear_LMDPL
constant Tile_X49Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000011111111101010100000000000000000111111110000000000000000101010100000000001010101000000000000000000000000000000000000000000000000010101010101010100000000101010101111111111111111000000000000000010101010101010100000000000000000";
--X50Y21, linear_LMDPL
constant Tile_X50Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000001010101010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X51Y21, nonlinear_LMDPL
constant Tile_X51Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000001111111100000000010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000001010101001010101000100010001000100000000101010100011001100110011000000000000000000000000000000000100010001000100";
--X52Y21, linear_LMDPL
constant Tile_X52Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101111111110000000000000000101010101010101001010101101010100000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000";
--X53Y21, linear_LMDPL
constant Tile_X53Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101111111110000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001010101010101010";
--X54Y21, nonlinear_LMDPL
constant Tile_X54Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111000000000000000010101010010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X55Y21, linear_LMDPL
constant Tile_X55Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000001010101010101010111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X56Y21, linear_LMDPL
constant Tile_X56Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000001010101000000001010101000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X57Y21, nonlinear_LMDPL
constant Tile_X57Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000101010100000000001010101000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X58Y21, linear_LMDPL
constant Tile_X58Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000001111111110101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000001010101000000000010001000100010011111111101010100000000000000000111111111111111101010101010101010000000000000000";
--X59Y21, linear_LMDPL
constant Tile_X59Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000101010100000000000100010001000100000000010101010100010001000100000000000000000000000000000000000010001000100010";
--X60Y21, nonlinear_LMDPL
constant Tile_X60Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000101010101010101010101010010001000100010000000000101010100000000000000000011001100110011000000000000000000000000000000000";
--X61Y21, linear_LMDPL
constant Tile_X61Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000010101011010101000000000101010100000000001010101101010100101010101010101010101011111111110101010000000001111111101010101000000001010101000000000000000001010101001010101000000000000000000000000010001000100010000000000010101010000000000000000000000000000000011001100110011000000000000000000";
--X62Y21, linear_LMDPL
constant Tile_X62Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000001010101000000000101010100101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000010101010101010111111111000000000000000000000000010101011010101000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X63Y21, nonlinear_LMDPL
constant Tile_X63Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000011001100110011000000000000000001000100010001000";
--X64Y21, linear_LMDPL
constant Tile_X64Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010110101010101010100000000001010101000000001010101000000000101010100000000000000000000000000101010100000000111111111010101001010101000000000000000000000000101010100000000000000000001000100010001000000000000000001100110011001100";
--X65Y21, linear_LMDPL
constant Tile_X65Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000101010100000000000000000111111110000000000000000101010100000000011111111000000000000000000000000000000000101010100000000000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X66Y21, nonlinear_LMDPL
constant Tile_X66Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000001100110011001110101010101010100000000000000000";
--X67Y21, linear_LMDPL
constant Tile_X67Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000111111110000000000000000101010101010101010101010000000000000000010101010000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000000101010101010101";
--X68Y21, linear_LMDPL
constant Tile_X68Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101011111111010001000100010000000000101010100000000000000000010001000100010010101010101010100000000000000000";
--X69Y21, nonlinear_LMDPL
constant Tile_X69Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000010101010000000000000000010101010101010100000000101010100010001000100010000000000000000010001000100010000000000000000000";
--X70Y21, linear_LMDPL
constant Tile_X70Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000";
--X71Y21, linear_LMDPL
constant Tile_X71Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000010101010000000000000000000000000101010100000000011111111000000000000000000000000101010101010101001010101010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X72Y21, nonlinear_LMDPL
constant Tile_X72Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X73Y21, linear_LMDPL
constant Tile_X73Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000001000100010001";
--X74Y21, linear_LMDPL
constant Tile_X74Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010101010101";
--X75Y21, nonlinear_LMDPL
constant Tile_X75Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010100101010101010101000100010001000100000000101010100011001100110011000000000000000000000000000000001010101010101010";
--X76Y21, linear_LMDPL
constant Tile_X76Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101111111110101010101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000101010100000000000000000100010001000100011001100110011000000000000000000";
--X77Y21, linear_LMDPL
constant Tile_X77Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000101010101010101";
--X78Y21, ctrl_to_sec
constant Tile_X78Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y21, combined_WDDL
constant Tile_X79Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000000000000001010000000000000000000000000000000001010000000000000000000000000101000000000000000000000000000000001000110101010000011110000000000000000101010100101010100000000";
--X80Y21, combined_WDDL
constant Tile_X80Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000101000000000000011110001000100001010101000000000000000000000111011101101110100000000";
--X81Y21, ctrl_IO
constant Tile_X81Y21_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y22, W_IO_custom
constant Tile_X0Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000001010101000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y22, linear_LMDPL
constant Tile_X1Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X2Y22, linear_LMDPL
constant Tile_X2Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001111111111111111";
--X3Y22, nonlinear_LMDPL
constant Tile_X3Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000010101010101010100010001000100010000000000000000";
--X4Y22, linear_LMDPL
constant Tile_X4Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000100000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X5Y22, linear_LMDPL
constant Tile_X5Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000111111110000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000";
--X6Y22, nonlinear_LMDPL
constant Tile_X6Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000010001000100010000010001000100010000000000000000";
--X7Y22, linear_LMDPL
constant Tile_X7Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X8Y22, linear_LMDPL
constant Tile_X8Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000010001000100010";
--X9Y22, nonlinear_LMDPL
constant Tile_X9Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000100010001000100";
--X10Y22, linear_LMDPL
constant Tile_X10Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010111111110000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X11Y22, linear_LMDPL
constant Tile_X11Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000111111111010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X12Y22, nonlinear_LMDPL
constant Tile_X12Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001000100010001000";
--X13Y22, linear_LMDPL
constant Tile_X13Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001111111100000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X14Y22, linear_LMDPL
constant Tile_X14Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101001010101010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X15Y22, nonlinear_LMDPL
constant Tile_X15Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101010101010101010100000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001";
--X16Y22, linear_LMDPL
constant Tile_X16Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101011111111000000000000000000000000010101011010101010101010010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X17Y22, linear_LMDPL
constant Tile_X17Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X18Y22, nonlinear_LMDPL
constant Tile_X18Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000011001100110011000000000000000000100010001000100";
--X19Y22, linear_LMDPL
constant Tile_X19Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010101010100000000011111111000000000000000000000000010101010000000000000000010001000100010000000000000000000010001000100010";
--X20Y22, linear_LMDPL
constant Tile_X20Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000010101010010101010101010111111111000000000000000000000000000000000000000010011001100110010000000000000000";
--X21Y22, nonlinear_LMDPL
constant Tile_X21Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001111111100000000010101010000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000011001100110011";
--X22Y22, linear_LMDPL
constant Tile_X22Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000101010101010101";
--X23Y22, linear_LMDPL
constant Tile_X23Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000110011001100110000000000000000001000100010001000";
--X24Y22, nonlinear_LMDPL
constant Tile_X24Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X25Y22, linear_LMDPL
constant Tile_X25Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X26Y22, linear_LMDPL
constant Tile_X26Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000001010101010101010";
--X27Y22, nonlinear_LMDPL
constant Tile_X27Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000001111111100000000101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X28Y22, linear_LMDPL
constant Tile_X28Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000001000100010001";
--X29Y22, linear_LMDPL
constant Tile_X29Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101011111111000100010001000100000000000000000100010001000100000000000000000000000000000000000001000100010001";
--X30Y22, nonlinear_LMDPL
constant Tile_X30Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X31Y22, linear_LMDPL
constant Tile_X31Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000000000000000000";
--X32Y22, linear_LMDPL
constant Tile_X32Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000001010101000100010001000100000000000000000000000000000000000000000000000000000000000000000101010101010101";
--X33Y22, nonlinear_LMDPL
constant Tile_X33Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X34Y22, linear_LMDPL
constant Tile_X34Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011111111110101010101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X35Y22, linear_LMDPL
constant Tile_X35Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000101010100000000000000000000000001010101000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000110011001100110";
--X36Y22, nonlinear_LMDPL
constant Tile_X36Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000100010001000100000000000000001110111011101110000000000000000000000000000000000010001000100010";
--X37Y22, linear_LMDPL
constant Tile_X37Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000010101010000000000000000010101010000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X38Y22, linear_LMDPL
constant Tile_X38Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010101010100101010111111111010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X39Y22, nonlinear_LMDPL
constant Tile_X39Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000111011101110111010101010101010100000000000000000";
--X40Y22, linear_LMDPL
constant Tile_X40Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010101010101000000000000000000101010100000000000000000000000000000000111111110101010110101010000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X41Y22, linear_LMDPL
constant Tile_X41Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000000100010001000100";
--X42Y22, nonlinear_LMDPL
constant Tile_X42Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000100110011001100100000000000000001100110011001100";
--X43Y22, linear_LMDPL
constant Tile_X43Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000000000011111111000000000000000010101010000000001010101000000000010101010101010100000000000000001010101010101010000000000000000011111111111111110000000000000000";
--X44Y22, linear_LMDPL
constant Tile_X44Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X45Y22, nonlinear_LMDPL
constant Tile_X45Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010100000000000000000000000001010101001010101000000000101010100000000000000000000000000000000101010100000000001010101010001000100010000000000101010100000000000000000101010101010101010101010101010100000000000000000";
--X46Y22, linear_LMDPL
constant Tile_X46Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100101010110101010000000000000000000000000000000000000000010101010000100010001000100000000101010101001100110011001000000000000000000000000000000001101110111011101";
--X47Y22, linear_LMDPL
constant Tile_X47Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001110101010101010100000000000000000";
--X48Y22, nonlinear_LMDPL
constant Tile_X48Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000010001000100010000000000000000001001100110011001";
--X49Y22, linear_LMDPL
constant Tile_X49Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X50Y22, linear_LMDPL
constant Tile_X50Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001000100010001000";
--X51Y22, nonlinear_LMDPL
constant Tile_X51Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000001010101011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101011011101110111011000000000000000000100010001000100000000000000000";
--X52Y22, linear_LMDPL
constant Tile_X52Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X53Y22, linear_LMDPL
constant Tile_X53Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000111111110101010100000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X54Y22, nonlinear_LMDPL
constant Tile_X54Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000101010101001100110011001000000000000000010001000100010000000000000000000";
--X55Y22, linear_LMDPL
constant Tile_X55Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101001010101101010100000000000000000101010100000000000000000101010100101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000000010001000100010";
--X56Y22, linear_LMDPL
constant Tile_X56Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000111111111010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X57Y22, nonlinear_LMDPL
constant Tile_X57Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000001010101000000001010101000000000010101010101010100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X58Y22, linear_LMDPL
constant Tile_X58Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X59Y22, linear_LMDPL
constant Tile_X59Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X60Y22, nonlinear_LMDPL
constant Tile_X60Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000010101011010101000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000000000000000000";
--X61Y22, linear_LMDPL
constant Tile_X61Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001010101010101010000000000000000010101010101010100000000000000000000000000000000000000000000000001010101101010100000000000000000000000001111111100000000010101011010101001010101000000000000000010101010111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X62Y22, linear_LMDPL
constant Tile_X62Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000001010101001010101000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000111111111111111111001100110011000000000000000000";
--X63Y22, nonlinear_LMDPL
constant Tile_X63Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011010101000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X64Y22, linear_LMDPL
constant Tile_X64Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000101010100101010101010101101010100000000010101010101010100101010110101010000000000000000000000000101010100000000000000000100010001000100000000000000000001001100110011001";
--X65Y22, linear_LMDPL
constant Tile_X65Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000010101010111111110000000000000000111111110000000000000000000000000000000000000000000100010001000100000000010101011000100010001000000000000000000000000000000000001010101010101010";
--X66Y22, nonlinear_LMDPL
constant Tile_X66Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000010101010101010100000000101010100011001100110011000000000000000000100010001000100000000000000000";
--X67Y22, linear_LMDPL
constant Tile_X67Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000101010101111111100000000000000000000000000000000000000001010101010101010000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X68Y22, linear_LMDPL
constant Tile_X68Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101011010101011111111010101010101010110101010000000001000100010001000000000000000000010101010101010100000000000000000";
--X69Y22, nonlinear_LMDPL
constant Tile_X69Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000010101010000000000000000000000000010001000100010000000000101010100000000000000000101010101010101000100010001000100000000000000000";
--X70Y22, linear_LMDPL
constant Tile_X70Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000001010101010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X71Y22, linear_LMDPL
constant Tile_X71Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000010101010101010101010101000000000010101010101010100000000101010101111111111111111000000000000000010001000100010000000000000000000";
--X72Y22, nonlinear_LMDPL
constant Tile_X72Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000010101010000100010001000100000000101010100010001000100010000000000000000000000000000000000010001000100010";
--X73Y22, linear_LMDPL
constant Tile_X73Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X74Y22, linear_LMDPL
constant Tile_X74Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001100110011001100";
--X75Y22, nonlinear_LMDPL
constant Tile_X75Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101011010101000000000000000000000000000000000101010100101010110101010010101010101010111111111101010100100010001000100000000000000000010111011101110110000000000000000";
--X76Y22, linear_LMDPL
constant Tile_X76Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010101111111100000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010110101010010001000100010000000000000000000000000000000000010001000100010001010101010101010000000000000000";
--X77Y22, linear_LMDPL
constant Tile_X77Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111101010100000000000000000010101010101010100000000101010101001100110011001000000000000000011001100110011000000000000000000";
--X78Y22, ctrl_to_sec
constant Tile_X78Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y22, combined_WDDL
constant Tile_X79Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000001010000000000000000000000000000000001111000000000000000000000000101001010000000000000000000010100001000110101010111110100000000000000000101010100000000000000000";
--X80Y22, combined_WDDL
constant Tile_X80Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000111100000000000000000000000000000000000000000000000000000000000011110000101000000000000000000001000100001010101000000000000000000000100110011110111000000000";
--X81Y22, ctrl_IO
constant Tile_X81Y22_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y23, W_IO_custom
constant Tile_X0Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000000001010101000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y23, linear_LMDPL
constant Tile_X1Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001110111011101110";
--X2Y23, linear_LMDPL
constant Tile_X2Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X3Y23, nonlinear_LMDPL
constant Tile_X3Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001001100110011001";
--X4Y23, linear_LMDPL
constant Tile_X4Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000001010101000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X5Y23, linear_LMDPL
constant Tile_X5Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X6Y23, nonlinear_LMDPL
constant Tile_X6Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001000100010001000";
--X7Y23, linear_LMDPL
constant Tile_X7Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000101010100000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X8Y23, linear_LMDPL
constant Tile_X8Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000010101010010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X9Y23, nonlinear_LMDPL
constant Tile_X9Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X10Y23, linear_LMDPL
constant Tile_X10Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X11Y23, linear_LMDPL
constant Tile_X11Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X12Y23, nonlinear_LMDPL
constant Tile_X12Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111110101010101010100000000000000000000000001010101010101010101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000001000100010001000000000000000001110111011101110";
--X13Y23, linear_LMDPL
constant Tile_X13Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101001010101000100010001000100000000000000000100010001000100000000000000000000000000000000000110011001100110";
--X14Y23, linear_LMDPL
constant Tile_X14Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101011111111101010100000000010101010000000000101010100000000000000000000000001010101000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X15Y23, nonlinear_LMDPL
constant Tile_X15Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101010101010101010100000000000000000000000001111111110101010101010100000000010101010000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X16Y23, linear_LMDPL
constant Tile_X16Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000001010101001010101010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X17Y23, linear_LMDPL
constant Tile_X17Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000111111110000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X18Y23, nonlinear_LMDPL
constant Tile_X18Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X19Y23, linear_LMDPL
constant Tile_X19Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000010101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X20Y23, linear_LMDPL
constant Tile_X20Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X21Y23, nonlinear_LMDPL
constant Tile_X21Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010111111110000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000100010001000100";
--X22Y23, linear_LMDPL
constant Tile_X22Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000011001100110011000000000000000001101110111011101";
--X23Y23, linear_LMDPL
constant Tile_X23Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000010101010010001000100010010101010000000000000000000000000001000100010001000000000000000000000000000000000";
--X24Y23, nonlinear_LMDPL
constant Tile_X24Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000011001100110011000000000000000001110111011101110";
--X25Y23, linear_LMDPL
constant Tile_X25Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000110111011101110100000000000000000111011101110111";
--X26Y23, linear_LMDPL
constant Tile_X26Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X27Y23, nonlinear_LMDPL
constant Tile_X27Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X28Y23, linear_LMDPL
constant Tile_X28Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X29Y23, linear_LMDPL
constant Tile_X29Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000011111111000000000000000000000000101010100000000010101010010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X30Y23, nonlinear_LMDPL
constant Tile_X30Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010101010101010110101010101010100000000000000000";
--X31Y23, linear_LMDPL
constant Tile_X31Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X32Y23, linear_LMDPL
constant Tile_X32Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X33Y23, nonlinear_LMDPL
constant Tile_X33Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010111111111000000000000000000000000000000000000000000000000010001000100010000000000000000000110011001100110";
--X34Y23, linear_LMDPL
constant Tile_X34Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111111111100000000000000001100110011001100";
--X35Y23, linear_LMDPL
constant Tile_X35Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101000000000010101010000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X36Y23, nonlinear_LMDPL
constant Tile_X36Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000001000100010001";
--X37Y23, linear_LMDPL
constant Tile_X37Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000010101010000000000000000010101010000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100";
--X38Y23, linear_LMDPL
constant Tile_X38Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000010101010000100010001000100000000101010101001100110011001000000000000000000000000000000001010101010101010";
--X39Y23, nonlinear_LMDPL
constant Tile_X39Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000101110111011101100000000000000000001000100010001";
--X40Y23, linear_LMDPL
constant Tile_X40Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000101010101010101001010101000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010100101010101010101010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X41Y23, linear_LMDPL
constant Tile_X41Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000000010001000100010";
--X42Y23, nonlinear_LMDPL
constant Tile_X42Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000101010100000000001010101000000000000000000000000000000000000000010101010000100010001000100000000101010100110011001100110000000000000000000000000000000000011001100110011";
--X43Y23, linear_LMDPL
constant Tile_X43Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111010101011010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X44Y23, linear_LMDPL
constant Tile_X44Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000011011101110111010000000000000000";
--X45Y23, nonlinear_LMDPL
constant Tile_X45Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000111111111010101000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000010001000100010010011001100110010000000000000000";
--X46Y23, linear_LMDPL
constant Tile_X46Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000101010101010101010101010000000000000000000000000000000000000000011111111010101010101010101010101000000001101110111011101000000000000000010101010101010100000000000000000";
--X47Y23, linear_LMDPL
constant Tile_X47Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X48Y23, nonlinear_LMDPL
constant Tile_X48Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000101010100000000000000000000000011111111101010100000000000000000010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X49Y23, linear_LMDPL
constant Tile_X49Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000010101011111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X50Y23, linear_LMDPL
constant Tile_X50Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001111111100000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001110111011101110";
--X51Y23, nonlinear_LMDPL
constant Tile_X51Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X52Y23, linear_LMDPL
constant Tile_X52Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000010101010010101010000000000000000101010101010101000000000101010100000000001010101000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100010001000100011111111111111110000000000000000";
--X53Y23, linear_LMDPL
constant Tile_X53Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X54Y23, nonlinear_LMDPL
constant Tile_X54Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110101010100000000010101010101010100000000000000001101110111011101000000000000000011001100110011000000000000000000";
--X55Y23, linear_LMDPL
constant Tile_X55Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010101010101000000000000100010001000111111111000000000101010101010101000000000000000000000000000000001111111111111111";
--X56Y23, linear_LMDPL
constant Tile_X56Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000010101010000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000010101010101010100101010100000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X57Y23, nonlinear_LMDPL
constant Tile_X57Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000010101010000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000100010001000100";
--X58Y23, linear_LMDPL
constant Tile_X58Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001010101011111111101010100000000000000000000000000000000010101010000000001010101000000000010101010101010100000000101010101100110011001100000000000000000000100010001000100000000000000000";
--X59Y23, linear_LMDPL
constant Tile_X59Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000101010100101010100000000000000000000000000000000000000001010101000000000000100010001000100000000101010100101010101010101000000000000000000000000000000001000100010001000";
--X60Y23, nonlinear_LMDPL
constant Tile_X60Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100101010101010101000000000000000000000000000000001010101000000000010101011010101000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y23, linear_LMDPL
constant Tile_X61Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000101010100101010110101010111111110000000010101010000000000000000000000000000000000101010110101010000000001010101010101010000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001000100010001000";
--X62Y23, linear_LMDPL
constant Tile_X62Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101001010101000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101001010101000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X63Y23, nonlinear_LMDPL
constant Tile_X63Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000101010101110111011101110000000000000000000000000000000000100010001000100";
--X64Y23, linear_LMDPL
constant Tile_X64Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000000000000000000010101010111111110000000001010101000000001111111100000000101010100101010100000000000000000101010110101010000000000000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000001000100010001000";
--X65Y23, linear_LMDPL
constant Tile_X65Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X66Y23, nonlinear_LMDPL
constant Tile_X66Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000001100110011001101010101010101010000000000000000";
--X67Y23, linear_LMDPL
constant Tile_X67Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101011111111000000001111111100000000000000001010101000000000000000000000000000000000101010100000000000000000101010101010101010101010000000000000000010101010000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X68Y23, linear_LMDPL
constant Tile_X68Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000010101010000000000000000010101010000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000011101110111011101010101010101010000000000000000";
--X69Y23, nonlinear_LMDPL
constant Tile_X69Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000111111111010101000000000010101010101010100000000101010100011001100110011000000000000000010001000100010000000000000000000";
--X70Y23, linear_LMDPL
constant Tile_X70Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000101010100000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100101010100000000010101010101010100000000000000001101110111011101000000000000000011001100110011000000000000000000";
--X71Y23, linear_LMDPL
constant Tile_X71Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X72Y23, nonlinear_LMDPL
constant Tile_X72Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X73Y23, linear_LMDPL
constant Tile_X73Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000001010101010101010101010100000000101010100010001000100010000000000000000000000000000000000000000000000000";
--X74Y23, linear_LMDPL
constant Tile_X74Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010101010101011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001000100010001000";
--X75Y23, nonlinear_LMDPL
constant Tile_X75Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101001010101010101010101010100000000101010100011001100110011000000000000000010101010101010100000000000000000";
--X76Y23, linear_LMDPL
constant Tile_X76Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000111111111010101010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000011001100110011";
--X77Y23, linear_LMDPL
constant Tile_X77Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001100110011001100000000000000000011011101110111010000000000000000";
--X78Y23, ctrl_to_sec
constant Tile_X78Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y23, combined_WDDL
constant Tile_X79Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000001010000000000000000000000000000000000000000000000000000000000000101010100000000000000000000010100000000010101010101010100000000000000000100010000000000011001100";
--X80Y23, combined_WDDL
constant Tile_X80Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000010100000101000000000000000000001000100001010101000000000000000000000000000001000100000000000";
--X81Y23, ctrl_IO
constant Tile_X81Y23_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y24, W_IO_custom
constant Tile_X0Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y24, linear_LMDPL
constant Tile_X1Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X2Y24, linear_LMDPL
constant Tile_X2Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001011101110111011";
--X3Y24, nonlinear_LMDPL
constant Tile_X3Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000000000000000000";
--X4Y24, linear_LMDPL
constant Tile_X4Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100010011001100110010000000000000000";
--X5Y24, linear_LMDPL
constant Tile_X5Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001001100110011001";
--X6Y24, nonlinear_LMDPL
constant Tile_X6Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000100010001000100";
--X7Y24, linear_LMDPL
constant Tile_X7Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110101010100000000101010100000000000000000111111111010101000000000101010100000000010101010000000000000000000000000010101010000000010101010010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X8Y24, linear_LMDPL
constant Tile_X8Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101111111110101010000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X9Y24, nonlinear_LMDPL
constant Tile_X9Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X10Y24, linear_LMDPL
constant Tile_X10Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X11Y24, linear_LMDPL
constant Tile_X11Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000001000100010001";
--X12Y24, nonlinear_LMDPL
constant Tile_X12Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X13Y24, linear_LMDPL
constant Tile_X13Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000111111111010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X14Y24, linear_LMDPL
constant Tile_X14Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010000100010001000100000000000000000110011001100110000000000000000000000000000000001110111011101110";
--X15Y24, nonlinear_LMDPL
constant Tile_X15Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X16Y24, linear_LMDPL
constant Tile_X16Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000001010101010101010000000000000000000000000000000001010101011111111010101010101010100000000000000001010101010101010000000000000000000110011001100110000000000000000";
--X17Y24, linear_LMDPL
constant Tile_X17Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000010101011010101010101010010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X18Y24, nonlinear_LMDPL
constant Tile_X18Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X19Y24, linear_LMDPL
constant Tile_X19Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000101010101101110111011101000000000000000010101010101010100000000000000000";
--X20Y24, linear_LMDPL
constant Tile_X20Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X21Y24, nonlinear_LMDPL
constant Tile_X21Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010000000000101010100000000000000000000000000000000111111110000000000000000010101010101010100000000101010101100110011001100000000000000000000010001000100010000000000000000";
--X22Y24, linear_LMDPL
constant Tile_X22Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000101010101010101010101010000000000000000000100010001000100000000000000000";
--X23Y24, linear_LMDPL
constant Tile_X23Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000101010100000000000000000001000100010001000000000000000000011001100110011";
--X24Y24, nonlinear_LMDPL
constant Tile_X24Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X25Y24, linear_LMDPL
constant Tile_X25Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000111011101110111000000000000000001011101110111011";
--X26Y24, linear_LMDPL
constant Tile_X26Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000000000000000000000000000000000000110011001100110000000000000000";
--X27Y24, nonlinear_LMDPL
constant Tile_X27Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000001110111011101110";
--X28Y24, linear_LMDPL
constant Tile_X28Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000011101110111011100000000000000000000000000000000";
--X29Y24, linear_LMDPL
constant Tile_X29Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000000100010001000100";
--X30Y24, nonlinear_LMDPL
constant Tile_X30Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X31Y24, linear_LMDPL
constant Tile_X31Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000010001000100010000000000000000000000000000000000001000100010001";
--X32Y24, linear_LMDPL
constant Tile_X32Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000010001000100010";
--X33Y24, nonlinear_LMDPL
constant Tile_X33Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X34Y24, linear_LMDPL
constant Tile_X34Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010110101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X35Y24, linear_LMDPL
constant Tile_X35Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000011111111101010100000000000000000000000000000000010101010000100010001000101010101000000000010001000100010000000000000000000000000000000001001100110011001";
--X36Y24, nonlinear_LMDPL
constant Tile_X36Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000000110011001100110000000000000000000000000000000000011001100110011";
--X37Y24, linear_LMDPL
constant Tile_X37Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000111111110000000000000000000000001111111110101010010101010000000010101010000000000000000000000000101010100000000010101010010101010101010100000000000000001010101010101010000000000000000001010101010101010000000000000000";
--X38Y24, linear_LMDPL
constant Tile_X38Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000010101010000000000000000010101010010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X39Y24, nonlinear_LMDPL
constant Tile_X39Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000001010101010101010000100010001000100000000101010100110011001100110000000000000000000000000000000000001000100010001";
--X40Y24, linear_LMDPL
constant Tile_X40Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X41Y24, linear_LMDPL
constant Tile_X41Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000001111111100000000000000000101010100000000101010100000000010101010000000000000000011111111101010100000000000000000010001000100010000000000101010100000000000000000001000100010001000100010001000100000000000000000";
--X42Y24, nonlinear_LMDPL
constant Tile_X42Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000001010101001010101000000000000000000000000000000000101010100000000101010100000000010101010000000000000000000000000000000000000000001010101010001000100010000000000101010100000000000000000110011001100110001110111011101110000000000000000";
--X43Y24, linear_LMDPL
constant Tile_X43Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000001010101101010100000000000000000010101010101010100000000000000001010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001100110011001100";
--X44Y24, linear_LMDPL
constant Tile_X44Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000000000000101010100000000000000000000000000000000001010101101010100000000000000000010101010000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X45Y24, nonlinear_LMDPL
constant Tile_X45Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101001100110011001000000000000000011001100110011000000000000000000";
--X46Y24, linear_LMDPL
constant Tile_X46Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111101010101010101000000000000000000101010101010101000000000000000001010101101010100000000000000000101010100000000000000000101010100000000010101010000000000000000000000000000000000101010110101010010001000100010000000000101010100000000000000000110111011101110111001100110011000000000000000000";
--X47Y24, linear_LMDPL
constant Tile_X47Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000000000000000000000";
--X48Y24, nonlinear_LMDPL
constant Tile_X48Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000010001000100010000000000101010100000000000000000000000000000000000010001000100010000000000000000";
--X49Y24, linear_LMDPL
constant Tile_X49Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011111111100000000000000001111111100000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101001010101010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X50Y24, linear_LMDPL
constant Tile_X50Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001010101000000000000000011111111000000000000000010101010000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X51Y24, nonlinear_LMDPL
constant Tile_X51Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111010101010000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000100010001000100000000000000001110111011101110000000000000000000000000000000001100110011001100";
--X52Y24, linear_LMDPL
constant Tile_X52Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100101010100000000000000000000000010101010111111111010101000000000010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X53Y24, linear_LMDPL
constant Tile_X53Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000010101010000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X54Y24, nonlinear_LMDPL
constant Tile_X54Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001110111011101110000000000000000010101010101010100000000000000000";
--X55Y24, linear_LMDPL
constant Tile_X55Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X56Y24, linear_LMDPL
constant Tile_X56Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000001111111101010101101010100000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000001010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X57Y24, nonlinear_LMDPL
constant Tile_X57Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010000000001010101000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000101010101010101";
--X58Y24, linear_LMDPL
constant Tile_X58Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000101010100000000010101010010101010000000000000000000000001010101000000000010101010000000000000000101010100000000000000000111111110000000000000000000100010001000110101010000000000101010101010101000000000000000000000000000000001000100010001000";
--X59Y24, linear_LMDPL
constant Tile_X59Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X60Y24, nonlinear_LMDPL
constant Tile_X60Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111101010101000000000101010110101010000000000000000000000000000000001010101000000000010101010101010100000000000000000000000000000000101010101010101000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000010001000100010";
--X61Y24, linear_LMDPL
constant Tile_X61Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000101010110101010101010100000000000000000101010101111111100000000010101011010101010101010000000000000000010101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X62Y24, linear_LMDPL
constant Tile_X62Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000000000001111111100000000010101010000000000000000000000001111111100000000101010100101010100000000000000000000000000000000101010101010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X63Y24, nonlinear_LMDPL
constant Tile_X63Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101010001000100010000000000101010100000000000000000011001100110011001000100010001000000000000000000";
--X64Y24, linear_LMDPL
constant Tile_X64Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000010101010101010100000000000000000000000000000000000000000101010101010101010101010000000000000000010101010000000000101010110101010000100010001000100000000101010100100010001000100000000000000000000000000000000000011001100110011";
--X65Y24, linear_LMDPL
constant Tile_X65Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000111111111010101000000000101010100000000000000000000000000000000011111111000000000101010100000000000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100";
--X66Y24, nonlinear_LMDPL
constant Tile_X66Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y24, linear_LMDPL
constant Tile_X67Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101111111100000000101010100000000000000000000000001010101010101010000000000000000011111111000000000000000000000000010101010101010110101010010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X68Y24, linear_LMDPL
constant Tile_X68Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000101010101010101000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010101010101010101010010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X69Y24, nonlinear_LMDPL
constant Tile_X69Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101001010101101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100101010110101010010001000100010000000000101010100000000000000000101110111011101110001000100010000000000000000000";
--X70Y24, linear_LMDPL
constant Tile_X70Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000001010101011111111000000000000000000000000010101010101010100000000010001000100010000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X71Y24, linear_LMDPL
constant Tile_X71Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010001000100010000000000000000000";
--X72Y24, nonlinear_LMDPL
constant Tile_X72Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000101010100000000000000000000000000000000010011001100110010000000000000000";
--X73Y24, linear_LMDPL
constant Tile_X73Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X74Y24, linear_LMDPL
constant Tile_X74Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000101010110101010010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X75Y24, nonlinear_LMDPL
constant Tile_X75Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000000101010101010101";
--X76Y24, linear_LMDPL
constant Tile_X76Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000111111111010101010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X77Y24, linear_LMDPL
constant Tile_X77Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010111111110000000000000000010101010101010100000000101010101101110111011101000000000000000010111011101110110000000000000000";
--X78Y24, ctrl_to_sec
constant Tile_X78Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y24, combined_WDDL
constant Tile_X79Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011110000000000000101000000000000000000000000101010100000000000001010000010100001000110101010101010100000000000000000110011000000000000000000";
--X80Y24, combined_WDDL
constant Tile_X80Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000111100000000000000000000000000000000000000000000000000000000000010100000101000000000000000000001000100001010101000001111000000000000010001001110111000000000";
--X81Y24, ctrl_IO
constant Tile_X81Y24_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y25, W_IO_custom
constant Tile_X0Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y25, linear_LMDPL
constant Tile_X1Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010010101010000000000000000101010101010101000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000110011001100110";
--X2Y25, linear_LMDPL
constant Tile_X2Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000111111110000000000000000000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001110111011101110";
--X3Y25, nonlinear_LMDPL
constant Tile_X3Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000111111111001100110011001000000000000000000010001000100010000000000000000";
--X4Y25, linear_LMDPL
constant Tile_X4Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000100110011001100100110011001100110000000000000000";
--X5Y25, linear_LMDPL
constant Tile_X5Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000010101010101010101111111100000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001110111011101110";
--X6Y25, nonlinear_LMDPL
constant Tile_X6Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001010101010101010000000000000000";
--X7Y25, linear_LMDPL
constant Tile_X7Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010101010100000000010101010000000000000000000000000010101010000000010101010010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X8Y25, linear_LMDPL
constant Tile_X8Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000000000001010101000000000111111110000000000000000000000001010101010101010000000001010101010101010010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X9Y25, nonlinear_LMDPL
constant Tile_X9Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X10Y25, linear_LMDPL
constant Tile_X10Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000110011001100110000000000000000";
--X11Y25, linear_LMDPL
constant Tile_X11Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X12Y25, nonlinear_LMDPL
constant Tile_X12Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000010101010000000011111111000000001010101010101010000000000000000000000000010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X13Y25, linear_LMDPL
constant Tile_X13Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000001111111110101010000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000010101011010101010101010010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X14Y25, linear_LMDPL
constant Tile_X14Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101010101010010101010101010100000000000000001010101010101010000000000000000001010101010101010000000000000000";
--X15Y25, nonlinear_LMDPL
constant Tile_X15Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000010101010101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100110011001100100000000000000001111111111111111";
--X16Y25, linear_LMDPL
constant Tile_X16Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X17Y25, linear_LMDPL
constant Tile_X17Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X18Y25, nonlinear_LMDPL
constant Tile_X18Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X19Y25, linear_LMDPL
constant Tile_X19Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001111111111111111000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X20Y25, linear_LMDPL
constant Tile_X20Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000001111111100000000000000000000000010101010010001000100010000000000000000000000000000000000101110111011101111111111111111110000000000000000";
--X21Y25, nonlinear_LMDPL
constant Tile_X21Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X22Y25, linear_LMDPL
constant Tile_X22Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000101010100000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001100110011001110101010101010100000000000000000";
--X23Y25, linear_LMDPL
constant Tile_X23Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000100010001000100000000010101010010001000100010000000000000000000000000000000001010101010101010";
--X24Y25, nonlinear_LMDPL
constant Tile_X24Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010001000100010000000000101010100000000000000000010001000100010010101010101010100000000000000000";
--X25Y25, linear_LMDPL
constant Tile_X25Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X26Y25, linear_LMDPL
constant Tile_X26Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X27Y25, nonlinear_LMDPL
constant Tile_X27Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000011111111010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X28Y25, linear_LMDPL
constant Tile_X28Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111101010101010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X29Y25, linear_LMDPL
constant Tile_X29Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001100110011001100";
--X30Y25, nonlinear_LMDPL
constant Tile_X30Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X31Y25, linear_LMDPL
constant Tile_X31Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000111111110000000010101010000000000000000011111111000000000000000000000000101110111011101100000000000000000000000000000000";
--X32Y25, linear_LMDPL
constant Tile_X32Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101011111111010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X33Y25, nonlinear_LMDPL
constant Tile_X33Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000101010101010101";
--X34Y25, linear_LMDPL
constant Tile_X34Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100010001000100011011101110111010000000000000000";
--X35Y25, linear_LMDPL
constant Tile_X35Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000001010101010101010000000000000000";
--X36Y25, nonlinear_LMDPL
constant Tile_X36Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y25, linear_LMDPL
constant Tile_X37Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X38Y25, linear_LMDPL
constant Tile_X38Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100000000000000000000000000000000000000000000000000010001000100010";
--X39Y25, nonlinear_LMDPL
constant Tile_X39Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000000011001100110011000000000000000000000000000000000001000100010001";
--X40Y25, linear_LMDPL
constant Tile_X40Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000101010100000000011111111010001000100010011111111000000000000000000000000000100010001000100000000000000000000000000000000";
--X41Y25, linear_LMDPL
constant Tile_X41Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000010101010000000000000000000000000101010100000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001100110011001100";
--X42Y25, nonlinear_LMDPL
constant Tile_X42Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101111111100000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000000010001000100010000000000000000";
--X43Y25, linear_LMDPL
constant Tile_X43Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101110111011101110110000000000000000";
--X44Y25, linear_LMDPL
constant Tile_X44Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X45Y25, nonlinear_LMDPL
constant Tile_X45Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000000100010001000100000000010101010110011001100110000000000000000000000000000000000000000000000000";
--X46Y25, linear_LMDPL
constant Tile_X46Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000111111110000000000000000000000000000000000000000111111111010101010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X47Y25, linear_LMDPL
constant Tile_X47Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X48Y25, nonlinear_LMDPL
constant Tile_X48Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111111010101000000000010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X49Y25, linear_LMDPL
constant Tile_X49Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X50Y25, linear_LMDPL
constant Tile_X50Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000010101010000000001111111100000000000000000000000000000000010101010101010111111111000000000100010001000100000000000000000000100010001000100000000000000000";
--X51Y25, nonlinear_LMDPL
constant Tile_X51Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000001010101000000000000000000000000011111111101010100101010100000000010101010000000000000000000000000101010101010101101010100000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000001110111011101110000000000000000000100010001000100000000000000000";
--X52Y25, linear_LMDPL
constant Tile_X52Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000001110111011101110000000000000000";
--X53Y25, linear_LMDPL
constant Tile_X53Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101001010101000000000101010100000000000000000000000000000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000101010101010101";
--X54Y25, nonlinear_LMDPL
constant Tile_X54Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100101010100000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101011010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X55Y25, linear_LMDPL
constant Tile_X55Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000001010101000000000101010100000000010101010101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X56Y25, linear_LMDPL
constant Tile_X56Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000001010101010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010101010100000000000000000000000010101010000000001010101010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000010001000100010";
--X57Y25, nonlinear_LMDPL
constant Tile_X57Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000101010101110111011101110000000000000000000000000000000000100010001000100";
--X58Y25, linear_LMDPL
constant Tile_X58Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000101010100000000000000000000000000000000010101010101010100000000001010101010001000100010000000000101010100000000000000000000100010001000101110111011101110000000000000000";
--X59Y25, linear_LMDPL
constant Tile_X59Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000101010100000000000100010001000100000000101010100000000000000000000000000000000000000000000000000101010101010101";
--X60Y25, nonlinear_LMDPL
constant Tile_X60Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y25, linear_LMDPL
constant Tile_X61Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000101010110101010101010101111111101010101000000001111111100000000010101011010101010101010000000000101010110101010000000000101010100000000000000000000000000000000101010100000000000000000001000100010001000000000000000001101110111011101";
--X62Y25, linear_LMDPL
constant Tile_X62Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000101010100101010100000000101010100000000000000000101010100000000000000000000000000000000000000000010101010000000000000000110011001100110000000000000000000110011001100110";
--X63Y25, nonlinear_LMDPL
constant Tile_X63Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101011010101001010101000100010001000100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X64Y25, linear_LMDPL
constant Tile_X64Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101011010101000000000101010100000000000000000000000000000000011111111000000001010101011111111101010100000000010101010000000000000000000000000101010100101010110101010101010100101010110101010000000000101010100000000000000000000000000000000101010100000000000000000010001000100010000000000000000000010001000100010";
--X65Y25, linear_LMDPL
constant Tile_X65Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X66Y25, nonlinear_LMDPL
constant Tile_X66Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101011010101001010101000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X67Y25, linear_LMDPL
constant Tile_X67Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101111111100000000111111110000000000000000101010101010101010101010000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000001000100010001000000000000000000000000000000000";
--X68Y25, linear_LMDPL
constant Tile_X68Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000111111111010101010101010000100010001000110101010010101011000100010001000000000000000000000000000000000000100010001000100";
--X69Y25, nonlinear_LMDPL
constant Tile_X69Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000011111111000000000000000000000000000000001010101010101010000100010001000100000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X70Y25, linear_LMDPL
constant Tile_X70Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010011111111000000000000000000000000010101010101010110001000100010000000000000000000";
--X71Y25, linear_LMDPL
constant Tile_X71Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X72Y25, nonlinear_LMDPL
constant Tile_X72Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000100010001000100000000000000000000100010001000100";
--X73Y25, linear_LMDPL
constant Tile_X73Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000101010101010101000000000000000000000000101010101111111110101010000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X74Y25, linear_LMDPL
constant Tile_X74Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000111111110000000010101010000000001010101000000000000000000101010110101010000000000000000000000000000000000000000010101010000100010001000100000000010101011011101110111011000000000000000000000000000000000001000100010001";
--X75Y25, nonlinear_LMDPL
constant Tile_X75Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101010101010010101010101010100000000101010100011001100110011000000000000000011111111111111110000000000000000";
--X76Y25, linear_LMDPL
constant Tile_X76Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010100000000010101010010101010101010100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X77Y25, linear_LMDPL
constant Tile_X77Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010101010101010111001100110011000000000000000000";
--X78Y25, ctrl_to_sec
constant Tile_X78Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y25, combined_WDDL
constant Tile_X79Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001111000000000000000000000000000000000000000000000000101010100000000000001010000010100001000110101010101010100000000000000000110111010101010100000000";
--X80Y25, combined_WDDL
constant Tile_X80Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000000000000000001111000000000000000010100000101000000000000000000001000100000000101011111010000000000000011001101110111000000000";
--X81Y25, ctrl_IO
constant Tile_X81Y25_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y26, W_IO_custom
constant Tile_X0Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y26, linear_LMDPL
constant Tile_X1Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X2Y26, linear_LMDPL
constant Tile_X2Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101011101110111011100000000000000000";
--X3Y26, nonlinear_LMDPL
constant Tile_X3Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000010001000100010";
--X4Y26, linear_LMDPL
constant Tile_X4Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X5Y26, linear_LMDPL
constant Tile_X5Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X6Y26, nonlinear_LMDPL
constant Tile_X6Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X7Y26, linear_LMDPL
constant Tile_X7Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000111111110000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001110111011101110";
--X8Y26, linear_LMDPL
constant Tile_X8Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000101010100000000101010100000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000110011001100110010111011101110110000000000000000";
--X9Y26, nonlinear_LMDPL
constant Tile_X9Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X10Y26, linear_LMDPL
constant Tile_X10Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X11Y26, linear_LMDPL
constant Tile_X11Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X12Y26, nonlinear_LMDPL
constant Tile_X12Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X13Y26, linear_LMDPL
constant Tile_X13Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X14Y26, linear_LMDPL
constant Tile_X14Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000101010101010101001010101000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X15Y26, nonlinear_LMDPL
constant Tile_X15Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X16Y26, linear_LMDPL
constant Tile_X16Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101010101010010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X17Y26, linear_LMDPL
constant Tile_X17Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010101010101010100000000000000001011101110111011000000000000000010011001100110010000000000000000";
--X18Y26, nonlinear_LMDPL
constant Tile_X18Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010111111111000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X19Y26, linear_LMDPL
constant Tile_X19Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000101010101000100010001000000000000000000001000100010001000000000000000000";
--X20Y26, linear_LMDPL
constant Tile_X20Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X21Y26, nonlinear_LMDPL
constant Tile_X21Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000101010100001000100010001000000000000000000000000000000000000000000000000";
--X22Y26, linear_LMDPL
constant Tile_X22Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000101010100000000001010101000100010001000100000000101010101100110011001100000000000000000000000000000000000011001100110011";
--X23Y26, linear_LMDPL
constant Tile_X23Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000011111111010101010101010100000000000000001111111111111111000000000000000011101110111011100000000000000000";
--X24Y26, nonlinear_LMDPL
constant Tile_X24Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X25Y26, linear_LMDPL
constant Tile_X25Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000011001100110011";
--X26Y26, linear_LMDPL
constant Tile_X26Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X27Y26, nonlinear_LMDPL
constant Tile_X27Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X28Y26, linear_LMDPL
constant Tile_X28Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010101010101000000000010001000100010000000000000000000000000000000000001000100010001001010101010101010000000000000000";
--X29Y26, linear_LMDPL
constant Tile_X29Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X30Y26, nonlinear_LMDPL
constant Tile_X30Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X31Y26, linear_LMDPL
constant Tile_X31Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X32Y26, linear_LMDPL
constant Tile_X32Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000011111111000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000111011101110111010101010101010100000000000000000";
--X33Y26, nonlinear_LMDPL
constant Tile_X33Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X34Y26, linear_LMDPL
constant Tile_X34Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000111111110000000000000000000000000000000010101010101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101";
--X35Y26, linear_LMDPL
constant Tile_X35Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000011111111000000000000000011111111000000000000000010101010010101010101010100000000000000000111011101110111000000000000000001010101010101010000000000000000";
--X36Y26, nonlinear_LMDPL
constant Tile_X36Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y26, linear_LMDPL
constant Tile_X37Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000001010101010001000100010000000000000000000000000000000000111111111111111110001000100010000000000000000000";
--X38Y26, linear_LMDPL
constant Tile_X38Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101011111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100111011101110111010000000000000000";
--X39Y26, nonlinear_LMDPL
constant Tile_X39Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X40Y26, linear_LMDPL
constant Tile_X40Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010101010101000000000000000001010101000000000101010100000000000000000000000000000000101010100000000000000000000000000000000011111111101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001000100010001000";
--X41Y26, linear_LMDPL
constant Tile_X41Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100000000010101010101010100000000000000000000000000000000001010101010101010101010100000000101010100010001000100010000000000000000011001100110011000000000000000000";
--X42Y26, nonlinear_LMDPL
constant Tile_X42Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X43Y26, linear_LMDPL
constant Tile_X43Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000010101010000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X44Y26, linear_LMDPL
constant Tile_X44Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X45Y26, nonlinear_LMDPL
constant Tile_X45Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000011111111000100010001000100000000101010100010001000100010000000000000000000000000000000001001100110011001";
--X46Y26, linear_LMDPL
constant Tile_X46Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011010101000000000000000000000000000000000000000000000000001010101010101011111111100000000101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000100010001000110101010101010101010101010101010000000000000000000000000000000000000000000000000";
--X47Y26, linear_LMDPL
constant Tile_X47Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010110101010000000000000000000000000101010100101010111111111000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X48Y26, nonlinear_LMDPL
constant Tile_X48Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X49Y26, linear_LMDPL
constant Tile_X49Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000001111111100000000000000000000000000000000101010100000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X50Y26, linear_LMDPL
constant Tile_X50Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000011111111010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X51Y26, nonlinear_LMDPL
constant Tile_X51Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X52Y26, linear_LMDPL
constant Tile_X52Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000101010100000000010101010010101010000000000000000000000000000000001010101101010100101010101010101000000000000000000000000000000000101010100000000010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X53Y26, linear_LMDPL
constant Tile_X53Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000101010101010101000000000000000000000000000000001010101000000000000000001010101011111111000000000000000000000000000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X54Y26, nonlinear_LMDPL
constant Tile_X54Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X55Y26, linear_LMDPL
constant Tile_X55Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000010101010111111110000000000000000000000000101010100000000010101010101010100000000000000001111111111111111000000000000000000100010001000100000000000000000";
--X56Y26, linear_LMDPL
constant Tile_X56Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101011111111111111110000000010101010000000001010101010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001101110111011101";
--X57Y26, nonlinear_LMDPL
constant Tile_X57Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000101010101010101000000000000000000000000010101010000000001010101000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X58Y26, linear_LMDPL
constant Tile_X58Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001001100110011001";
--X59Y26, linear_LMDPL
constant Tile_X59Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001010101010101010000000000000000101010100000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111111010101001010101010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X60Y26, nonlinear_LMDPL
constant Tile_X60Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000101010100000000000100010001000100000000101010101110111011101110000000000000000000000000000000000010001000100010";
--X61Y26, linear_LMDPL
constant Tile_X61Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101011111111101010100000000000000000000000000101010100000000101010100000000001010101101010100000000000000000000000000000000000000000101010100000000010101010000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000111011101110111011001100110011000000000000000000";
--X62Y26, linear_LMDPL
constant Tile_X62Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000001010101000000000000000000000000000000000101010101010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001111111111111111";
--X63Y26, nonlinear_LMDPL
constant Tile_X63Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000001010101010101010101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X64Y26, linear_LMDPL
constant Tile_X64Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000000000000101010101111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000101010100000000010101010000000000000000010101010111111111010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000001100110011001100";
--X65Y26, linear_LMDPL
constant Tile_X65Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001111111111111111";
--X66Y26, nonlinear_LMDPL
constant Tile_X66Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y26, linear_LMDPL
constant Tile_X67Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010110101010000000000000000000000000111111111010101010101010000000000000000000000000010101010000000000000000101110111011101100000000000000000101010101010101";
--X68Y26, linear_LMDPL
constant Tile_X68Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X69Y26, nonlinear_LMDPL
constant Tile_X69Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101011010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000001010101000000000010101010101010100000000010101010000000000000000000000000000000010101010101010100000000000000000";
--X70Y26, linear_LMDPL
constant Tile_X70Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X71Y26, linear_LMDPL
constant Tile_X71Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111111010101000000000000000000000000010101010101010100000000000000000000100010001000100000000010101010011001100110011000000000000000000000000000000000010001000100010";
--X72Y26, nonlinear_LMDPL
constant Tile_X72Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X73Y26, linear_LMDPL
constant Tile_X73Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111111010101000000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101011111111010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X74Y26, linear_LMDPL
constant Tile_X74Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000000000000101010100000000010101010010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X75Y26, nonlinear_LMDPL
constant Tile_X75Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000101010100100010001000100000000000000000001010101010101010000000000000000";
--X76Y26, linear_LMDPL
constant Tile_X76Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111000000001111111110101010000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X77Y26, linear_LMDPL
constant Tile_X77Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X78Y26, ctrl_to_sec
constant Tile_X78Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y26, combined_WDDL
constant Tile_X79Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001011111000010100101010110101010101010100000000001010101000000000100010000000000";
--X80Y26, combined_WDDL
constant Tile_X80Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000001111101000000000000010100000101000000000000000000100010000000000101010101010000011011101000000000000000011101110";
--X81Y26, ctrl_IO
constant Tile_X81Y26_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y27, W_IO_custom
constant Tile_X0Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y27, linear_LMDPL
constant Tile_X1Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000001011101110111011";
--X2Y27, linear_LMDPL
constant Tile_X2Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010101010000000000000000000000001111111100000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000001100110011001100000000000000000";
--X3Y27, nonlinear_LMDPL
constant Tile_X3Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001000100010001000";
--X4Y27, linear_LMDPL
constant Tile_X4Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000010101010101010100000000000000000011001100110011000000000000000001100110011001100000000000000000";
--X5Y27, linear_LMDPL
constant Tile_X5Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000010101010010101010101010100000000000000000001000100010001000000000000000001000100010001000000000000000000";
--X6Y27, nonlinear_LMDPL
constant Tile_X6Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000001111111101010101000000000000000001010101000000000000000001010101000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001011101110111011";
--X7Y27, linear_LMDPL
constant Tile_X7Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010010101010000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X8Y27, linear_LMDPL
constant Tile_X8Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000101010101111111100000000101010100000000000000000000000000101010110101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X9Y27, nonlinear_LMDPL
constant Tile_X9Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101001010101111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X10Y27, linear_LMDPL
constant Tile_X10Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010101010000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000001010101001010101000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000010101010100010001000100000000000000000000010001000100010000000000000000";
--X11Y27, linear_LMDPL
constant Tile_X11Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111110101010101010100000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X12Y27, nonlinear_LMDPL
constant Tile_X12Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000001111111100000000101010100000000010101010000000001010101000000000000000000000000000000000000000000101010110101010101010100000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X13Y27, linear_LMDPL
constant Tile_X13Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X14Y27, linear_LMDPL
constant Tile_X14Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X15Y27, nonlinear_LMDPL
constant Tile_X15Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000101010100000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X16Y27, linear_LMDPL
constant Tile_X16Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X17Y27, linear_LMDPL
constant Tile_X17Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000010101011010101010101010010101010101010100000000000000000010001000100010000000000000000010011001100110010000000000000000";
--X18Y27, nonlinear_LMDPL
constant Tile_X18Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000001000100010001";
--X19Y27, linear_LMDPL
constant Tile_X19Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X20Y27, linear_LMDPL
constant Tile_X20Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001111111110101010000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X21Y27, nonlinear_LMDPL
constant Tile_X21Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X22Y27, linear_LMDPL
constant Tile_X22Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000110011001100110000110011001100110000000000000000";
--X23Y27, linear_LMDPL
constant Tile_X23Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000000000000000000010101010101010100000000000000000";
--X24Y27, nonlinear_LMDPL
constant Tile_X24Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000001000100010001000000000000000001100110011001100";
--X25Y27, linear_LMDPL
constant Tile_X25Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X26Y27, linear_LMDPL
constant Tile_X26Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X27Y27, nonlinear_LMDPL
constant Tile_X27Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000101010100000000010101010101010100000000000000000011001100110011000000000000000010011001100110010000000000000000";
--X28Y27, linear_LMDPL
constant Tile_X28Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X29Y27, linear_LMDPL
constant Tile_X29Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101011111111111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X30Y27, nonlinear_LMDPL
constant Tile_X30Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X31Y27, linear_LMDPL
constant Tile_X31Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000110011001100110";
--X32Y27, linear_LMDPL
constant Tile_X32Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000111011101110111";
--X33Y27, nonlinear_LMDPL
constant Tile_X33Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X34Y27, linear_LMDPL
constant Tile_X34Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000001010101000000000000000000000000000000000000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000000110011001100110";
--X35Y27, linear_LMDPL
constant Tile_X35Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000010101010101010110101010000000000000000000000000000000000000000010101010101010100000000000000000";
--X36Y27, nonlinear_LMDPL
constant Tile_X36Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X37Y27, linear_LMDPL
constant Tile_X37Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X38Y27, linear_LMDPL
constant Tile_X38Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010001000100010000000000101010100000000000000000011001100110011000000000000000000000000000000000";
--X39Y27, nonlinear_LMDPL
constant Tile_X39Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y27, linear_LMDPL
constant Tile_X40Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001111111111111111";
--X41Y27, linear_LMDPL
constant Tile_X41Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100101010101010101000000000000000000000000000000000000000000000000";
--X42Y27, nonlinear_LMDPL
constant Tile_X42Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100011001100110011000000000000000000000000000000000001000100010001";
--X43Y27, linear_LMDPL
constant Tile_X43Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000001010101011111111010001000100010000000000000000000000000000000000000100010001000101010101010101010000000000000000";
--X44Y27, linear_LMDPL
constant Tile_X44Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X45Y27, nonlinear_LMDPL
constant Tile_X45Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000010101010000000001010101000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000101010100000000000100010001000100000000101010101010101010101010000000000000000000000000000000001010101010101010";
--X46Y27, linear_LMDPL
constant Tile_X46Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010101111111101010101000000000000000000000000000000000000000000000000101010100101010100000000000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X47Y27, linear_LMDPL
constant Tile_X47Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000010101010101010100000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000101010101010101";
--X48Y27, nonlinear_LMDPL
constant Tile_X48Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000100010001000100";
--X49Y27, linear_LMDPL
constant Tile_X49Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X50Y27, linear_LMDPL
constant Tile_X50Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000111111110000000000000000000000000000000010101010000000000000000010101010101010100101010110101010010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X51Y27, nonlinear_LMDPL
constant Tile_X51Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X52Y27, linear_LMDPL
constant Tile_X52Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000101010100101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X53Y27, linear_LMDPL
constant Tile_X53Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011";
--X54Y27, nonlinear_LMDPL
constant Tile_X54Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X55Y27, linear_LMDPL
constant Tile_X55Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000010101010000000010101010000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X56Y27, linear_LMDPL
constant Tile_X56Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000101010100101010110101010000000000000000010101010000000001010101010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X57Y27, nonlinear_LMDPL
constant Tile_X57Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000000000000000000001010101000000001111111110101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000110111011101110100000000000000001010101010101010";
--X58Y27, linear_LMDPL
constant Tile_X58Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000001010101101010100101010101010101101010100000000010101010000000000000000000000000000100010001000110101010000000001100110011001100000000000000000000000000000000001000100010001000";
--X59Y27, linear_LMDPL
constant Tile_X59Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010101010101010101010000100010001000100000000101010100101010101010101000000000000000000000000000000000010001000100010";
--X60Y27, nonlinear_LMDPL
constant Tile_X60Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000010001000100010";
--X61Y27, linear_LMDPL
constant Tile_X61Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010101010100000000000000000101010100000000010101010000000000101010110101010111111111010101000000000000000000000000011111111101010100000000000000000001000100010001000000000000000001101110111011101";
--X62Y27, linear_LMDPL
constant Tile_X62Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000101010101010101000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001001100110011001";
--X63Y27, nonlinear_LMDPL
constant Tile_X63Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X64Y27, linear_LMDPL
constant Tile_X64Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001111111100000000101010100000000001010101000000000000000010101010010101011010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001100110011001100";
--X65Y27, linear_LMDPL
constant Tile_X65Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000110111011101110100000000000000000111011101110111";
--X66Y27, nonlinear_LMDPL
constant Tile_X66Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000010101011010101010101010010101010101010100000000101010101110111011101110000000000000000001010101010101010000000000000000";
--X67Y27, linear_LMDPL
constant Tile_X67Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000011111111101010100101010110101010000000000000000000000000000000001010101010101010010001000100010000000000010101010000000000000000010001000100010011001100110011000000000000000000";
--X68Y27, linear_LMDPL
constant Tile_X68Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000010101011000100010001000000000000000000000000000000000000000000000000000";
--X69Y27, nonlinear_LMDPL
constant Tile_X69Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X70Y27, linear_LMDPL
constant Tile_X70Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010001000100010011111111000000000000000000000000000000000000000011001100110011000000000000000000";
--X71Y27, linear_LMDPL
constant Tile_X71Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X72Y27, nonlinear_LMDPL
constant Tile_X72Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000101110111011101100000000000000000100010001000100";
--X73Y27, linear_LMDPL
constant Tile_X73Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000011111111000000001010101000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X74Y27, linear_LMDPL
constant Tile_X74Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000101010100000000000000001010101010101010000000000000000000000000101010100101010100000000010101010101010100000000000000001010101010101010000000000000000001010101010101010000000000000000";
--X75Y27, nonlinear_LMDPL
constant Tile_X75Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010101010101000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X76Y27, linear_LMDPL
constant Tile_X76Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111111111111101010100000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000001000100010001";
--X77Y27, linear_LMDPL
constant Tile_X77Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X78Y27, ctrl_to_sec
constant Tile_X78Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y27, combined_WDDL
constant Tile_X79Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000001111000000000000000000000000000000000000101000000000000000000000000010100101010110101010101010100000000010001000000000001111111100000000";
--X80Y27, combined_WDDL
constant Tile_X80Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000111100000000000000000000000000000000101010101010000000000000001100110000000011111111";
--X81Y27, ctrl_IO
constant Tile_X81Y27_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y28, W_IO_custom
constant Tile_X0Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y28, linear_LMDPL
constant Tile_X1Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X2Y28, linear_LMDPL
constant Tile_X2Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000001000100010001";
--X3Y28, nonlinear_LMDPL
constant Tile_X3Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000001000100010001000000000000000000";
--X4Y28, linear_LMDPL
constant Tile_X4Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010010101010000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X5Y28, linear_LMDPL
constant Tile_X5Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X6Y28, nonlinear_LMDPL
constant Tile_X6Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010110101010000000000000000000000000000000001111111110101010010101010000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001110111011101110";
--X7Y28, linear_LMDPL
constant Tile_X7Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000101010100000000000000000000000000000000010101010000000000000000010101010000000001111111100000000000000000000000010101010000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X8Y28, linear_LMDPL
constant Tile_X8Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001011101110111011";
--X9Y28, nonlinear_LMDPL
constant Tile_X9Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000101010100000000000000000000000001010101000000000101010101010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X10Y28, linear_LMDPL
constant Tile_X10Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X11Y28, linear_LMDPL
constant Tile_X11Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101001010101010101010000000001010101000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000110011001100110000110011001100110000000000000000";
--X12Y28, nonlinear_LMDPL
constant Tile_X12Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000011111111101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X13Y28, linear_LMDPL
constant Tile_X13Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000000000000000000001010101000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X14Y28, linear_LMDPL
constant Tile_X14Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000000110011001100110000000000000000010001000100010000000000000000000";
--X15Y28, nonlinear_LMDPL
constant Tile_X15Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000100010001000100";
--X16Y28, linear_LMDPL
constant Tile_X16Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000001010101000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X17Y28, linear_LMDPL
constant Tile_X17Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000001010101010101010010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X18Y28, nonlinear_LMDPL
constant Tile_X18Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y28, linear_LMDPL
constant Tile_X19Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000010111011101110110000000000000000";
--X20Y28, linear_LMDPL
constant Tile_X20Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001011101110111011000000000000000000000000000000000001000100010001";
--X21Y28, nonlinear_LMDPL
constant Tile_X21Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X22Y28, linear_LMDPL
constant Tile_X22Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X23Y28, linear_LMDPL
constant Tile_X23Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X24Y28, nonlinear_LMDPL
constant Tile_X24Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X25Y28, linear_LMDPL
constant Tile_X25Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101100110011001100000000000000000001000100010001000000000000000000";
--X26Y28, linear_LMDPL
constant Tile_X26Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000111111110100010001000100000000000000000010011001100110010000000000000000";
--X27Y28, nonlinear_LMDPL
constant Tile_X27Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001000100010001000";
--X28Y28, linear_LMDPL
constant Tile_X28Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101010101010101010100000000000000000111011101110111000000000000000011011101110111010000000000000000";
--X29Y28, linear_LMDPL
constant Tile_X29Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111111111111010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000011001100110011";
--X30Y28, nonlinear_LMDPL
constant Tile_X30Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001001100110011001";
--X31Y28, linear_LMDPL
constant Tile_X31Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000000101010101010101000000000000000011111111111111110000000000000000";
--X32Y28, linear_LMDPL
constant Tile_X32Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000010101010000000000101010100000000101010100000000000000000000100010001000100000000111111110100010001000100000000000000000000000000000000000001000100010001";
--X33Y28, nonlinear_LMDPL
constant Tile_X33Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000001000100010001";
--X34Y28, linear_LMDPL
constant Tile_X34Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000101010100000000111111110000000011111111111111110000000010101010010101010000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X35Y28, linear_LMDPL
constant Tile_X35Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000111111110000000000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X36Y28, nonlinear_LMDPL
constant Tile_X36Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y28, linear_LMDPL
constant Tile_X37Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X38Y28, linear_LMDPL
constant Tile_X38Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X39Y28, nonlinear_LMDPL
constant Tile_X39Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000010101011110111011101110000000000000000000000000000000000011001100110011";
--X40Y28, linear_LMDPL
constant Tile_X40Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000010101010101010100000000001010101000000000000000000000000000000000000000000000000001100110011001100000000000000000110011001100110";
--X41Y28, linear_LMDPL
constant Tile_X41Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000101010100000000010101010000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X42Y28, nonlinear_LMDPL
constant Tile_X42Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X43Y28, linear_LMDPL
constant Tile_X43Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000010101010000000010101010000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X44Y28, linear_LMDPL
constant Tile_X44Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111101010101101010100000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000010101010100010001000100000000000000000000000000000000001100110011001100";
--X45Y28, nonlinear_LMDPL
constant Tile_X45Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000001100110011001100";
--X46Y28, linear_LMDPL
constant Tile_X46Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000111111110000000010101010101010101010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000011101110111011100000000000000001110111011101110";
--X47Y28, linear_LMDPL
constant Tile_X47Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101011010101000000000010101010101010100000000010101011100110011001100000000000000000010001000100010000000000000000000";
--X48Y28, nonlinear_LMDPL
constant Tile_X48Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000010101010101010100000000101010101011101110111011000000000000000000000000000000000000000000000000";
--X49Y28, linear_LMDPL
constant Tile_X49Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X50Y28, linear_LMDPL
constant Tile_X50Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000101010101010101011111111111111110000000000000000";
--X51Y28, nonlinear_LMDPL
constant Tile_X51Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000000000001010101011111111000100010001000100000000000000000110011001100110000000000000000000000000000000000001000100010001";
--X52Y28, linear_LMDPL
constant Tile_X52Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000000000000000000";
--X53Y28, linear_LMDPL
constant Tile_X53Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010101010101000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000110111011101110111001100110011000000000000000000";
--X54Y28, nonlinear_LMDPL
constant Tile_X54Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100101010111111111000000000000000000000000000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000001100110011001100";
--X55Y28, linear_LMDPL
constant Tile_X55Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000101010101111111100000000000000001010101000000000111111110000000010101010101010100000000000000000010101010101010100000000000100010001000100000000000000001010101010101010000000000000000000000000000000001101110111011101";
--X56Y28, linear_LMDPL
constant Tile_X56Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010111111110000000000000000111111110000000000000000101010101010101010101010000000000000000010101010000000001010101010101010010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X57Y28, nonlinear_LMDPL
constant Tile_X57Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000010101010000000000000000000000001010101001010101000000000000000001010101010101010000000000000000000000000101010100000000111111110101010100000000000000000000000001010101000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000100010001000100";
--X58Y28, linear_LMDPL
constant Tile_X58Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000000010001000100010";
--X59Y28, linear_LMDPL
constant Tile_X59Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010101010101000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000111111111010101000000000101010100000000001010101000000000000000000000000111111111010101010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X60Y28, nonlinear_LMDPL
constant Tile_X60Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000010001000100010";
--X61Y28, linear_LMDPL
constant Tile_X61Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000010101010000000000000000111111110000000000000000111111110101010100000000000000001010101000000000101010100101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X62Y28, linear_LMDPL
constant Tile_X62Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000001010101000000000111111110000000011111111101010100000000000000000010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X63Y28, nonlinear_LMDPL
constant Tile_X63Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001010101010101010";
--X64Y28, linear_LMDPL
constant Tile_X64Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000101010100000000000000000101010101010101000000000010001000100010000000000101010100000000000000000000000000000000010001000100010000000000000000000";
--X65Y28, linear_LMDPL
constant Tile_X65Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000011111111000000000101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X66Y28, nonlinear_LMDPL
constant Tile_X66Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000001100110011001100000000000000000000000000000000";
--X67Y28, linear_LMDPL
constant Tile_X67Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000010101010000000000000000000000000101010101010101010101010000000000000000011111111000000001010101001010101010001000100010000000000010101010000000000000000110011001100110010101010101010100000000000000000";
--X68Y28, linear_LMDPL
constant Tile_X68Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010010101010101010110101010000000000100010001000100000000000000000000100010001000100000000000000000";
--X69Y28, nonlinear_LMDPL
constant Tile_X69Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y28, linear_LMDPL
constant Tile_X70Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001111111111111111000000000000000000000000000000000000000000000000";
--X71Y28, linear_LMDPL
constant Tile_X71Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000001010101010101010";
--X72Y28, nonlinear_LMDPL
constant Tile_X72Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000000000000101010101010101000000000010101010101010100000000101010100000000000000000000000000000000010101010101010100000000000000000";
--X73Y28, linear_LMDPL
constant Tile_X73Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000001010101001010101000000000000000000000000101010100000000000000000001100110011001100000000000000000000000000000000";
--X74Y28, linear_LMDPL
constant Tile_X74Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X75Y28, nonlinear_LMDPL
constant Tile_X75Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000001010101000000000000000000000000101010101010101000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000001000100010001";
--X76Y28, linear_LMDPL
constant Tile_X76Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001101110111011101000000000000000010001000100010000000000000000000";
--X77Y28, linear_LMDPL
constant Tile_X77Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X78Y28, ctrl_to_sec
constant Tile_X78Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y28, combined_WDDL
constant Tile_X79Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000011110101010110101010101010100000111101000100000000000011001100000000";
--X80Y28, combined_WDDL
constant Tile_X80Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000101010100000111110101111000000000000000000000101010100000000101010101010000011001100000000001011101100000000";
--X81Y28, ctrl_IO
constant Tile_X81Y28_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y29, W_IO_custom
constant Tile_X0Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y29, linear_LMDPL
constant Tile_X1Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001100110011001100";
--X2Y29, linear_LMDPL
constant Tile_X2Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X3Y29, nonlinear_LMDPL
constant Tile_X3Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y29, linear_LMDPL
constant Tile_X4Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101000000000101010100000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001001100110011001";
--X5Y29, linear_LMDPL
constant Tile_X5Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101001010101101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X6Y29, nonlinear_LMDPL
constant Tile_X6Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010000000010101010000000001111111100000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000000010001000100010000000000000000";
--X7Y29, linear_LMDPL
constant Tile_X7Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010101010100000000101010100000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000001111111110101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X8Y29, linear_LMDPL
constant Tile_X8Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000001010101101010100000000000000000000000000000000010101010000000000000000000000000010101010101010100000000010101010011001100110011000000000000000000100010001000100000000000000000";
--X9Y29, nonlinear_LMDPL
constant Tile_X9Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101011111111100000000101010100000000000000000000000001010101000000000101010101010101000000000000000000000000000000000101010100000000000000000000100010001000100000000010101010001000100010001000000000000000000000000000000000100010001000100";
--X10Y29, linear_LMDPL
constant Tile_X10Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000010101010101010100000000010101010000000000101010110101010101010100000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X11Y29, linear_LMDPL
constant Tile_X11Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111111010101000000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X12Y29, nonlinear_LMDPL
constant Tile_X12Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000010101010101010100000000011111111010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X13Y29, linear_LMDPL
constant Tile_X13Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X14Y29, linear_LMDPL
constant Tile_X14Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X15Y29, nonlinear_LMDPL
constant Tile_X15Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X16Y29, linear_LMDPL
constant Tile_X16Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000001010101010101010010101010101010100000000000000000100010001000100000000000000000000010001000100010000000000000000";
--X17Y29, linear_LMDPL
constant Tile_X17Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X18Y29, nonlinear_LMDPL
constant Tile_X18Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y29, linear_LMDPL
constant Tile_X19Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X20Y29, linear_LMDPL
constant Tile_X20Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X21Y29, nonlinear_LMDPL
constant Tile_X21Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X22Y29, linear_LMDPL
constant Tile_X22Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000111111110000000010101010000000000000000000000000111111110000000000000000000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000110011001100110";
--X23Y29, linear_LMDPL
constant Tile_X23Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X24Y29, nonlinear_LMDPL
constant Tile_X24Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000000110011001100110";
--X25Y29, linear_LMDPL
constant Tile_X25Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X26Y29, linear_LMDPL
constant Tile_X26Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000001010101000100010001000100000000000000001011101110111011000000000000000000000000000000001010101010101010";
--X27Y29, nonlinear_LMDPL
constant Tile_X27Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000110011001100110";
--X28Y29, linear_LMDPL
constant Tile_X28Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X29Y29, linear_LMDPL
constant Tile_X29Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X30Y29, nonlinear_LMDPL
constant Tile_X30Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X31Y29, linear_LMDPL
constant Tile_X31Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X32Y29, linear_LMDPL
constant Tile_X32Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X33Y29, nonlinear_LMDPL
constant Tile_X33Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y29, linear_LMDPL
constant Tile_X34Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010101010000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X35Y29, linear_LMDPL
constant Tile_X35Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001010101000000000101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X36Y29, nonlinear_LMDPL
constant Tile_X36Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X37Y29, linear_LMDPL
constant Tile_X37Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010111111110000000000000000101010101111111110101010010001000100010000000000000000000000000000000000010001000100010010011001100110010000000000000000";
--X38Y29, linear_LMDPL
constant Tile_X38Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000001010101001010101000100010001000100000000101010101010101010101010000000000000000000000000000000001010101010101010";
--X39Y29, nonlinear_LMDPL
constant Tile_X39Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y29, linear_LMDPL
constant Tile_X40Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X41Y29, linear_LMDPL
constant Tile_X41Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111101010101101010100000000000000000101010100000000000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010001000100010000000000000000000";
--X42Y29, nonlinear_LMDPL
constant Tile_X42Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111010101010000000000000000000000000000000000000000101010100000000000000000101010100000000001010101000000000000000000000000010101011010101010101010000100010001000100000000101010100011001100110011000000000000000000000000000000000110011001100110";
--X43Y29, linear_LMDPL
constant Tile_X43Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010101111111100000000000000001010101000000000000000000101010100000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000101010101010101001010101010101010000000000000000";
--X44Y29, linear_LMDPL
constant Tile_X44Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101001010101000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X45Y29, nonlinear_LMDPL
constant Tile_X45Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000101010100011001100110011000000000000000010001000100010000000000000000000";
--X46Y29, linear_LMDPL
constant Tile_X46Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101001010101010101010000000000000000000000000000000000000000010101010000000000000000111111110000000000000000101010101010101000000000000000000101010100000000000000000000000000000000000000000101010101010101010001000100010000000000000000000000000000000000001000100010001011111111111111110000000000000000";
--X47Y29, linear_LMDPL
constant Tile_X47Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000101010100000000011111111000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X48Y29, nonlinear_LMDPL
constant Tile_X48Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001100110011001100110011001100110000000000000000";
--X49Y29, linear_LMDPL
constant Tile_X49Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010101010101000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000011111111010101010101010101010101000100010001000100000000000000001100110011001100000000000000000000000000000000001011101110111011";
--X50Y29, linear_LMDPL
constant Tile_X50Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010010101010000000000000000101010100000000000000000000000000000000010101010000000001010101000000000101010100000000000000000000000000000000000000000101010100101010111111111000000000000000000000000000000001010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X51Y29, nonlinear_LMDPL
constant Tile_X51Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010000000000000000000000000000000000000000001010101101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000000000000000000";
--X52Y29, linear_LMDPL
constant Tile_X52Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000010001000100010";
--X53Y29, linear_LMDPL
constant Tile_X53Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010101010101010101011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X54Y29, nonlinear_LMDPL
constant Tile_X54Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111010101001010101000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000111011101110111";
--X55Y29, linear_LMDPL
constant Tile_X55Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000101010100000000010101010101010100000000000000000000000001010101000000000010101010101010101010101000000000000000000000000101010100101010100000000010001000100010000000000010101010000000000000000111111111111111110001000100010000000000000000000";
--X56Y29, linear_LMDPL
constant Tile_X56Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X57Y29, nonlinear_LMDPL
constant Tile_X57Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001010101000000000101010100000000011111111000000000000000000000000101010100101010101010101101010100000000010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000000000000100110011001100100000000000000000001000100010001";
--X58Y29, linear_LMDPL
constant Tile_X58Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000111111110000000000000000000000001111111100000000101010100101010100000000000000000000000010101010000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X59Y29, linear_LMDPL
constant Tile_X59Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010110101010000000000000000000000000111111111010101010101010010001000100010000000000101010100000000000000000101110111011101101010101010101010000000000000000";
--X60Y29, nonlinear_LMDPL
constant Tile_X60Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111010101001010101000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000110111011101110100000000000000000111011101110111";
--X61Y29, linear_LMDPL
constant Tile_X61Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001100110011001100";
--X62Y29, linear_LMDPL
constant Tile_X62Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000101010100101010100000000000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001101110111011101";
--X63Y29, nonlinear_LMDPL
constant Tile_X63Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101011010101000000000010101010101010100000000101010101110111011101110000000000000000000100010001000100000000000000000";
--X64Y29, linear_LMDPL
constant Tile_X64Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010101010101000000000010001000100010000000000101010100000000000000000110111011101110111011101110111010000000000000000";
--X65Y29, linear_LMDPL
constant Tile_X65Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000001010101000000000000000000000000000000000000000000000000010101010111111110000000000000000111111111010101000000000000000000000000001010101111111110000000000000000000000000101010101010101010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X66Y29, nonlinear_LMDPL
constant Tile_X66Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000001100110011001100000000000000001011101110111011";
--X67Y29, linear_LMDPL
constant Tile_X67Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000101010101111111100000000101010100000000000000000000000001010101000000000000000000000000010101010111111111010101000000000101010100101010110101010000000000000000000000000000000001010101001010101000000000000000000000000010101010000000000000000010001000100010000000000000000000010001000100010";
--X68Y29, linear_LMDPL
constant Tile_X68Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010010101010101010100000000000000000101010101010101000000000000000000100010001000100000000000000000";
--X69Y29, nonlinear_LMDPL
constant Tile_X69Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X70Y29, linear_LMDPL
constant Tile_X70Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000001010101010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X71Y29, linear_LMDPL
constant Tile_X71Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X72Y29, nonlinear_LMDPL
constant Tile_X72Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101001010101010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X73Y29, linear_LMDPL
constant Tile_X73Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000000000000011111111000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X74Y29, linear_LMDPL
constant Tile_X74Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X75Y29, nonlinear_LMDPL
constant Tile_X75Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010101010101010100000000101010101000100010001000000000000000000010111011101110110000000000000000";
--X76Y29, linear_LMDPL
constant Tile_X76Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X77Y29, linear_LMDPL
constant Tile_X77Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101010001000100010000000000010101010000000000000000001100110011001111001100110011000000000000000000";
--X78Y29, ctrl_to_sec
constant Tile_X78Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000101111100000000000000000000000000000000000000000000000000001111000000000000000000000000";
--X79Y29, combined_WDDL
constant Tile_X79Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000000000000000000000000000000000000000000000000000000000010100000000000001111101000000000000000000000000000000101010110100000101010100000000010101010000000000101010100000000";
--X80Y29, combined_WDDL
constant Tile_X80Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000101000000000000000010100000000000000000000000000001000100000000101010101010111100000000110111011001100100000000";
--X81Y29, ctrl_IO
constant Tile_X81Y29_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y30, W_IO_custom
constant Tile_X0Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y30, linear_LMDPL
constant Tile_X1Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X2Y30, linear_LMDPL
constant Tile_X2Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X3Y30, nonlinear_LMDPL
constant Tile_X3Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y30, linear_LMDPL
constant Tile_X4Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X5Y30, linear_LMDPL
constant Tile_X5Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010101010101010100010001000100010000000000000000";
--X6Y30, nonlinear_LMDPL
constant Tile_X6Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001010101000000000000000000101010100000000000100010001000100000000000000001000100010001000000000000000000000000000000000001001100110011001";
--X7Y30, linear_LMDPL
constant Tile_X7Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000001010101101010100000000010101010101010100000000000000000000000000101010110101010010101010000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X8Y30, linear_LMDPL
constant Tile_X8Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000101010100000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X9Y30, nonlinear_LMDPL
constant Tile_X9Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000001010101001010101010101011010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000000110011001100110000000000000000";
--X10Y30, linear_LMDPL
constant Tile_X10Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010111111110000000000000000000000000000000010101010010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X11Y30, linear_LMDPL
constant Tile_X11Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000010101010000000000000000000000000000000001010101000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X12Y30, nonlinear_LMDPL
constant Tile_X12Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X13Y30, linear_LMDPL
constant Tile_X13Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X14Y30, linear_LMDPL
constant Tile_X14Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X15Y30, nonlinear_LMDPL
constant Tile_X15Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X16Y30, linear_LMDPL
constant Tile_X16Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X17Y30, linear_LMDPL
constant Tile_X17Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X18Y30, nonlinear_LMDPL
constant Tile_X18Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y30, linear_LMDPL
constant Tile_X19Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000010101010010001000100010000000000101010100000000000000000100010001000100001000100010001000000000000000000";
--X20Y30, linear_LMDPL
constant Tile_X20Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000110011001100110";
--X21Y30, nonlinear_LMDPL
constant Tile_X21Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X22Y30, linear_LMDPL
constant Tile_X22Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000010101010101010110101010101010100000000000000000";
--X23Y30, linear_LMDPL
constant Tile_X23Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X24Y30, nonlinear_LMDPL
constant Tile_X24Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X25Y30, linear_LMDPL
constant Tile_X25Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100101010101010101000000000000000010111011101110110000000000000000";
--X26Y30, linear_LMDPL
constant Tile_X26Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001100110011001100000000000000000011101110111011100000000000000000";
--X27Y30, nonlinear_LMDPL
constant Tile_X27Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X28Y30, linear_LMDPL
constant Tile_X28Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011101110111011100100010001000100000000000000000";
--X29Y30, linear_LMDPL
constant Tile_X29Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000010001000100010000000000000000011011101110111010000000000000000";
--X30Y30, nonlinear_LMDPL
constant Tile_X30Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X31Y30, linear_LMDPL
constant Tile_X31Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000110011001100110";
--X32Y30, linear_LMDPL
constant Tile_X32Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X33Y30, nonlinear_LMDPL
constant Tile_X33Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y30, linear_LMDPL
constant Tile_X34Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X35Y30, linear_LMDPL
constant Tile_X35Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000101010101010101010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000";
--X36Y30, nonlinear_LMDPL
constant Tile_X36Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y30, linear_LMDPL
constant Tile_X37Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101010111011101110110000000000000000";
--X38Y30, linear_LMDPL
constant Tile_X38Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000010101011010101000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000111111110000000001010101010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X39Y30, nonlinear_LMDPL
constant Tile_X39Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000010101011110111011101110000000000000000000000000000000000101010101010101";
--X40Y30, linear_LMDPL
constant Tile_X40Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000111111110101010100000000111111110000000010101010000000000000000010101010010101010101010100000000000000000111011101110111000000000000000000110011001100110000000000000000";
--X41Y30, linear_LMDPL
constant Tile_X41Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000010101010000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011101110111011100100010001000100000000000000000";
--X42Y30, nonlinear_LMDPL
constant Tile_X42Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X43Y30, linear_LMDPL
constant Tile_X43Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000000000001010101000000000111111111010101011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111";
--X44Y30, linear_LMDPL
constant Tile_X44Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101011111111100000000000000000000000000000000000000000101010100000000101010101111111100000000101010100000000000000000010101011010101000000000101010100000000010101010101010100101010100000000010101010101010100000000101010100000000000000000000000000000000010001000100010000000000000000000";
--X45Y30, nonlinear_LMDPL
constant Tile_X45Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001010101010101010";
--X46Y30, linear_LMDPL
constant Tile_X46Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010101010101000000000000000000000000101010101111111101010101111111110000000000000000000000001111111100000000000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X47Y30, linear_LMDPL
constant Tile_X47Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111111010101011111111000000000000000000000000101010101010101000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001100110011001100";
--X48Y30, nonlinear_LMDPL
constant Tile_X48Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001110111011101110000000000000000000100010001000100000000000000000";
--X49Y30, linear_LMDPL
constant Tile_X49Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001010101010101010010001000100010001010101000000000000000000000000010001000100010011001100110011000000000000000000";
--X50Y30, linear_LMDPL
constant Tile_X50Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010101011010101000000000000000000000000000000000010101010000000000000000101010100000000000000000000000001111111100000000101010101010101000000000000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X51Y30, nonlinear_LMDPL
constant Tile_X51Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000110011001100110000000000000000011001100110011000000000000000000";
--X52Y30, linear_LMDPL
constant Tile_X52Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000001111111100000000000000000000000000000000000000001010101000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X53Y30, linear_LMDPL
constant Tile_X53Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000111111110101010110101010101010101010101010101010000000000000000001010101000000000101010100000000010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X54Y30, nonlinear_LMDPL
constant Tile_X54Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101101010100000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X55Y30, linear_LMDPL
constant Tile_X55Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000010101010010101010000000000000000101010101010101000000000000000001010101000000000000000000000000000000000111111110101010100000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X56Y30, linear_LMDPL
constant Tile_X56Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000001010101000000000000000010101010010101010000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000001010101010101010000100010001000100000000000000000101010101010101000000000000000000000000000000000100010001000100";
--X57Y30, nonlinear_LMDPL
constant Tile_X57Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000001111111100000000000000001010101000000000000000001010101010101010010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101011010101000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000100010001000100";
--X58Y30, linear_LMDPL
constant Tile_X58Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000001111111100000000000000000000000000000000111111110000000000000000000000001111111100000000101010100101010101010101101010100000000000000000000000001010101000000000000100010001000110101010000000001100110011001100000000000000000000000000000000000010001000100010";
--X59Y30, linear_LMDPL
constant Tile_X59Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101101010100101010100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000101010110101010000000000000000000000000101010100101010110101010000100010001000100000000000000000111011101110111000000000000000000000000000000000111011101110111";
--X60Y30, nonlinear_LMDPL
constant Tile_X60Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000001010101000000000101010100000000000100010001000100000000101010101110111011101110000000000000000000000000000000000100010001000100";
--X61Y30, linear_LMDPL
constant Tile_X61Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000101010100000000000000000000000001010101000000000000000000000000001010101000000001111111100000000000000000000000000000000010001000100010010101010000000000000000000000000010001000100010000100010001000100000000000000000";
--X62Y30, linear_LMDPL
constant Tile_X62Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000001111111100000000101010101111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000100010001000100000000000000001010101010101010";
--X63Y30, nonlinear_LMDPL
constant Tile_X63Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000011111111000000000000000000000000101010100101010100000000000100010001000100000000101010100110011001100110000000000000000000000000000000001001100110011001";
--X64Y30, linear_LMDPL
constant Tile_X64Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010101010101001010101000100010001000100000000101010101010101010101010000000000000000000000000000000001011101110111011";
--X65Y30, linear_LMDPL
constant Tile_X65Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000111111110000000001010101000000000000000010101010000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000111011101110111";
--X66Y30, nonlinear_LMDPL
constant Tile_X66Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y30, linear_LMDPL
constant Tile_X67Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000101010101010101001010101000000000000000010101010000000001010101010101010000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000";
--X68Y30, linear_LMDPL
constant Tile_X68Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010101010101010101010010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X69Y30, nonlinear_LMDPL
constant Tile_X69Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y30, linear_LMDPL
constant Tile_X70Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000011111111111111110000000000000000";
--X71Y30, linear_LMDPL
constant Tile_X71Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X72Y30, nonlinear_LMDPL
constant Tile_X72Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X73Y30, linear_LMDPL
constant Tile_X73Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010101101110111011101000000000000000010111011101110110000000000000000";
--X74Y30, linear_LMDPL
constant Tile_X74Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X75Y30, nonlinear_LMDPL
constant Tile_X75Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000101010101000100010001000000000000000000010101010101010100000000000000000";
--X76Y30, linear_LMDPL
constant Tile_X76Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X77Y30, linear_LMDPL
constant Tile_X77Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000010001000100010010111011101110110000000000000000";
--X78Y30, ctrl_to_sec
constant Tile_X78Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y30, combined_WDDL
constant Tile_X79Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000101001010000000000000000000000000101010111110000101010100000000000000000000000001111111100000000";
--X80Y30, combined_WDDL
constant Tile_X80Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000000000000000000000101000000000000000000000000000000000000000000000000000000000111100000000000011110000000000000101010100000000000010101010101010001000000000001101110100000000";
--X81Y30, ctrl_IO
constant Tile_X81Y30_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y31, W_IO_custom
constant Tile_X0Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y31, linear_LMDPL
constant Tile_X1Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X2Y31, linear_LMDPL
constant Tile_X2Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X3Y31, nonlinear_LMDPL
constant Tile_X3Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001101110111011101";
--X4Y31, linear_LMDPL
constant Tile_X4Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111101010101010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X5Y31, linear_LMDPL
constant Tile_X5Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001010101000000000010101010000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000101010101010101000000000000000010101010101010100000000000000000";
--X6Y31, nonlinear_LMDPL
constant Tile_X6Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X7Y31, linear_LMDPL
constant Tile_X7Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000001010101010101010000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000010101010100010001000100000000000000000010101010101010100000000000000000";
--X8Y31, linear_LMDPL
constant Tile_X8Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010101010101010111111111010101010000000000000000000000001111111100000000010001000100010000000000101010100000000000000000100010001000100011011101110111010000000000000000";
--X9Y31, nonlinear_LMDPL
constant Tile_X9Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000001010101000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100000000000000000001100110011001100000000000000000";
--X10Y31, linear_LMDPL
constant Tile_X10Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010101010100000000000000000101010100000000010101010111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001001100110011001";
--X11Y31, linear_LMDPL
constant Tile_X11Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001100110011001100";
--X12Y31, nonlinear_LMDPL
constant Tile_X12Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101001010101000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000001000100010001";
--X13Y31, linear_LMDPL
constant Tile_X13Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000001000100010001000000000000000000000000000000000101010101010101";
--X14Y31, linear_LMDPL
constant Tile_X14Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001110111011101110";
--X15Y31, nonlinear_LMDPL
constant Tile_X15Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X16Y31, linear_LMDPL
constant Tile_X16Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000010101010101010100000000000000000110011001100110000000000000000010011001100110010000000000000000";
--X17Y31, linear_LMDPL
constant Tile_X17Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X18Y31, nonlinear_LMDPL
constant Tile_X18Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y31, linear_LMDPL
constant Tile_X19Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000101010100000000011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101010101010101010100000000000000000";
--X20Y31, linear_LMDPL
constant Tile_X20Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001111111111111111";
--X21Y31, nonlinear_LMDPL
constant Tile_X21Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X22Y31, linear_LMDPL
constant Tile_X22Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000010001000100010011111111000000000000000000000000000000000000000001000100010001000000000000000000";
--X23Y31, linear_LMDPL
constant Tile_X23Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100";
--X24Y31, nonlinear_LMDPL
constant Tile_X24Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X25Y31, linear_LMDPL
constant Tile_X25Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X26Y31, linear_LMDPL
constant Tile_X26Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X27Y31, nonlinear_LMDPL
constant Tile_X27Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X28Y31, linear_LMDPL
constant Tile_X28Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X29Y31, linear_LMDPL
constant Tile_X29Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X30Y31, nonlinear_LMDPL
constant Tile_X30Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X31Y31, linear_LMDPL
constant Tile_X31Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X32Y31, linear_LMDPL
constant Tile_X32Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X33Y31, nonlinear_LMDPL
constant Tile_X33Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X34Y31, linear_LMDPL
constant Tile_X34Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X35Y31, linear_LMDPL
constant Tile_X35Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100101010111111111000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110010001000100010000000000000000000";
--X36Y31, nonlinear_LMDPL
constant Tile_X36Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X37Y31, linear_LMDPL
constant Tile_X37Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000010101010000000010101010000000000000000011111111101010101111111110101010010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X38Y31, linear_LMDPL
constant Tile_X38Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000111111111010101000000000000000000000000010101010000000001010101001010101000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X39Y31, nonlinear_LMDPL
constant Tile_X39Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000110011001100110000000000000000001010101010101010000000000000000";
--X40Y31, linear_LMDPL
constant Tile_X40Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X41Y31, linear_LMDPL
constant Tile_X41Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X42Y31, nonlinear_LMDPL
constant Tile_X42Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000001110111011101110000000000000000000100010001000100000000000000000";
--X43Y31, linear_LMDPL
constant Tile_X43Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000101010110101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X44Y31, linear_LMDPL
constant Tile_X44Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000101010100000000001010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001010101010101010";
--X45Y31, nonlinear_LMDPL
constant Tile_X45Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000010001000100010";
--X46Y31, linear_LMDPL
constant Tile_X46Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000111011101110111010101010101010100000000000000000";
--X47Y31, linear_LMDPL
constant Tile_X47Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000101010100000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010101010101001010101000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X48Y31, nonlinear_LMDPL
constant Tile_X48Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101010101010101010100000000000000000000000000000000000000000101010101010101001010101000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X49Y31, linear_LMDPL
constant Tile_X49Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X50Y31, linear_LMDPL
constant Tile_X50Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111010101011111111100000000000000000000000000000000000000000000000001010101010101011111111100000000000000000000000010101010101010101010101000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000110011001100110";
--X51Y31, nonlinear_LMDPL
constant Tile_X51Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101010101010000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000010101010101010100010001000100010000000000000000";
--X52Y31, linear_LMDPL
constant Tile_X52Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000100110011001100100000000000000000101010101010101";
--X53Y31, linear_LMDPL
constant Tile_X53Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X54Y31, nonlinear_LMDPL
constant Tile_X54Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000101010110101010000000000000000000000000111111111010101000000000000000000101010100000000000000000000000010101010000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010011001100110010000000000000000";
--X55Y31, linear_LMDPL
constant Tile_X55Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000000000000011111111000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000001010101000000000101010100000000000000000101010101010101000000000000100010001000100000000101010100000000000000000000000000000000000000000000000000101010101010101";
--X56Y31, linear_LMDPL
constant Tile_X56Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000101010100000000001010101101010100000000000000000000000000101010100000000101010100101010100000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X57Y31, nonlinear_LMDPL
constant Tile_X57Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000001010101000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000001001100110011001";
--X58Y31, linear_LMDPL
constant Tile_X58Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000001010101011111111000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101001010101000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000110011001100110000000000000000000101010101010101";
--X59Y31, linear_LMDPL
constant Tile_X59Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000010101010101010100000000010101010000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000110011001100110000000000000000000101010101010101";
--X60Y31, nonlinear_LMDPL
constant Tile_X60Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000001000100010001";
--X61Y31, linear_LMDPL
constant Tile_X61Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000001010101010001000100010000000000101010100000000000000000100110011001100110101010101010100000000000000000";
--X62Y31, linear_LMDPL
constant Tile_X62Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000101010100000000000000000101010101010101011111111000000000000000011111111000000000000000001010101000100010001000100000000101010100000000000000000000000000000000000000000000000001010101010101010";
--X63Y31, nonlinear_LMDPL
constant Tile_X63Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000101010100000000001010101000000000000000000000000111111111010101000000000000000000000000000000000101010100000000000000000001000100010001000000000000000001001100110011001";
--X64Y31, linear_LMDPL
constant Tile_X64Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110101010111111111000000000101010100000000111111110000000000000000101010101010101010101010000000000000000000000000101010100000000000000000110011001100110000000000000000001010101010101010";
--X65Y31, linear_LMDPL
constant Tile_X65Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101011111111000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100101010111111111010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X66Y31, nonlinear_LMDPL
constant Tile_X66Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010101010101010101010010101010101010100000000010101010110011001100110000000000000000001000100010001000000000000000000";
--X67Y31, linear_LMDPL
constant Tile_X67Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111101010100000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100000000000000000000000000000000000000000000000001010101010101010";
--X68Y31, linear_LMDPL
constant Tile_X68Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111101010101010101010101010000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000";
--X69Y31, nonlinear_LMDPL
constant Tile_X69Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y31, linear_LMDPL
constant Tile_X70Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X71Y31, linear_LMDPL
constant Tile_X71Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000101010100000000000000000000000000000000001010101010101010000000000000000";
--X72Y31, nonlinear_LMDPL
constant Tile_X72Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X73Y31, linear_LMDPL
constant Tile_X73Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000001011101110111011";
--X74Y31, linear_LMDPL
constant Tile_X74Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X75Y31, nonlinear_LMDPL
constant Tile_X75Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001001100110011001";
--X76Y31, linear_LMDPL
constant Tile_X76Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000100010001000100000000000000000000001000100010001";
--X77Y31, linear_LMDPL
constant Tile_X77Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X78Y31, ctrl_to_sec
constant Tile_X78Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000";
--X79Y31, combined_WDDL
constant Tile_X79Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010110100000111110100000010100000000000000001101110100000000";
--X80Y31, combined_WDDL
constant Tile_X80Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000111100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001000100000000000010101010000000000000100110011001100100000000";
--X81Y31, ctrl_IO
constant Tile_X81Y31_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y32, W_IO_custom
constant Tile_X0Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y32, linear_LMDPL
constant Tile_X1Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001111111111111111";
--X2Y32, linear_LMDPL
constant Tile_X2Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X3Y32, nonlinear_LMDPL
constant Tile_X3Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X4Y32, linear_LMDPL
constant Tile_X4Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X5Y32, linear_LMDPL
constant Tile_X5Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000111111110000000010101010010101010101010100000000000000000001000100010001000000000000000010001000100010000000000000000000";
--X6Y32, nonlinear_LMDPL
constant Tile_X6Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010111111110000000000000000000000001010101000000000000000000000000000000000000100010001000100000000010101011011101110111011000000000000000000000000000000001010101010101010";
--X7Y32, linear_LMDPL
constant Tile_X7Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000001111111100000000010101010101010100000000000000001001100110011001000000000000000000110011001100110000000000000000";
--X8Y32, linear_LMDPL
constant Tile_X8Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110101010100000000000000000000000000000000101010100000000001010101010101010000000000000000000000000101010101010101000000001010101010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111011101110111000000000000000001000100010001000";
--X9Y32, nonlinear_LMDPL
constant Tile_X9Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001011101110111011";
--X10Y32, linear_LMDPL
constant Tile_X10Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000011111111010101010000000000000000000000000000000001010101101010101010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X11Y32, linear_LMDPL
constant Tile_X11Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X12Y32, nonlinear_LMDPL
constant Tile_X12Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010";
--X13Y32, linear_LMDPL
constant Tile_X13Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X14Y32, linear_LMDPL
constant Tile_X14Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X15Y32, nonlinear_LMDPL
constant Tile_X15Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X16Y32, linear_LMDPL
constant Tile_X16Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000100010001000100";
--X17Y32, linear_LMDPL
constant Tile_X17Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X18Y32, nonlinear_LMDPL
constant Tile_X18Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X19Y32, linear_LMDPL
constant Tile_X19Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000010101010101010100000000010101010000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000010001000100010011011101110111010000000000000000";
--X20Y32, linear_LMDPL
constant Tile_X20Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001010101010101010";
--X21Y32, nonlinear_LMDPL
constant Tile_X21Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000000000000000000";
--X22Y32, linear_LMDPL
constant Tile_X22Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X23Y32, linear_LMDPL
constant Tile_X23Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X24Y32, nonlinear_LMDPL
constant Tile_X24Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000001000100010001000000000000000000000000000000001000100010001000";
--X25Y32, linear_LMDPL
constant Tile_X25Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010001000100010000000000101010100000000000000000001100110011001110101010101010100000000000000000";
--X26Y32, linear_LMDPL
constant Tile_X26Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000101010100000000001010101010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X27Y32, nonlinear_LMDPL
constant Tile_X27Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X28Y32, linear_LMDPL
constant Tile_X28Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X29Y32, linear_LMDPL
constant Tile_X29Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001110111011101110000000000000000";
--X30Y32, nonlinear_LMDPL
constant Tile_X30Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000101010101010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000101010101010101";
--X31Y32, linear_LMDPL
constant Tile_X31Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X32Y32, linear_LMDPL
constant Tile_X32Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X33Y32, nonlinear_LMDPL
constant Tile_X33Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X34Y32, linear_LMDPL
constant Tile_X34Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X35Y32, linear_LMDPL
constant Tile_X35Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X36Y32, nonlinear_LMDPL
constant Tile_X36Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000101010100000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000011001100110011";
--X37Y32, linear_LMDPL
constant Tile_X37Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000001010101010101010010001000100010000000000000000000000000000000000100010001000100011001100110011000000000000000000";
--X38Y32, linear_LMDPL
constant Tile_X38Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000010001000100010";
--X39Y32, nonlinear_LMDPL
constant Tile_X39Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001110111011101110000000000000000001010101010101010000000000000000";
--X40Y32, linear_LMDPL
constant Tile_X40Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X41Y32, linear_LMDPL
constant Tile_X41Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X42Y32, nonlinear_LMDPL
constant Tile_X42Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X43Y32, linear_LMDPL
constant Tile_X43Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010100000000000000000101010100000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X44Y32, linear_LMDPL
constant Tile_X44Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000101010101010101101010100000000000000000101010100000000000000000010101010000000011111111000000000000000010101010101010100000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000000101010101010101";
--X45Y32, nonlinear_LMDPL
constant Tile_X45Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000010101010000000000000000010101010101010100000000000000001110111011101110000000000000000000100010001000100000000000000000";
--X46Y32, linear_LMDPL
constant Tile_X46Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010101010101000000000010101010000000000000000000000000000000001010101000000001010101000000000010001000100010000000000000000000000000000000000010101010101010101010101010101010000000000000000";
--X47Y32, linear_LMDPL
constant Tile_X47Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000100010001000100000000000000000000000000000000000";
--X48Y32, nonlinear_LMDPL
constant Tile_X48Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010101010101000000000111111110000000000000000000000001010101001010101101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000001110111011101110";
--X49Y32, linear_LMDPL
constant Tile_X49Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X50Y32, linear_LMDPL
constant Tile_X50Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000001010101011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000001000100010001";
--X51Y32, nonlinear_LMDPL
constant Tile_X51Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000001010101000000001010101001010101000100010001000100000000000000001100110011001100000000000000000000000000000000001101110111011101";
--X52Y32, linear_LMDPL
constant Tile_X52Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010101010110101010000000000000000000000000010101010101010111111111000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X53Y32, linear_LMDPL
constant Tile_X53Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000101010100000000000000000111111110000000000000000000000000000000000000000101010101010101001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X54Y32, nonlinear_LMDPL
constant Tile_X54Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001010101000000000101010100101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X55Y32, linear_LMDPL
constant Tile_X55Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001111111101010101010101010000000000000000101010101010101000000000000000001010101000000000111111110000000000000000101010101010101000000000010001000100010000000000000000000000000000000000000100010001000101010101010101010000000000000000";
--X56Y32, linear_LMDPL
constant Tile_X56Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000001111111100000000010101010000000001010101000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X57Y32, nonlinear_LMDPL
constant Tile_X57Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010010101010101010101010101000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X58Y32, linear_LMDPL
constant Tile_X58Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000011001100110011000000000000000001101110111011101";
--X59Y32, linear_LMDPL
constant Tile_X59Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010110101010101010100000000010101010000000000000000000000000101010101010101011111111010001000100010000000000000000000000000000000000100110011001100110101010101010100000000000000000";
--X60Y32, nonlinear_LMDPL
constant Tile_X60Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X61Y32, linear_LMDPL
constant Tile_X61Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000001010101000000000010101010101010100000000000000000000000000000000111111110101010100000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X62Y32, linear_LMDPL
constant Tile_X62Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010101010101010101010101010100000000000000000000000000000000000000000101010101010101010101010111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001011101110111011";
--X63Y32, nonlinear_LMDPL
constant Tile_X63Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000010101010000000010101010000000000000000000000000010101011010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001000100010001000";
--X64Y32, linear_LMDPL
constant Tile_X64Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001111111100000000101010100000000000000000000000000101010100000000101010101010101000000000000000000000000010101010111111111010101010101010010001000100010000000000000000000000000000000000110011001100110001010101010101010000000000000000";
--X65Y32, linear_LMDPL
constant Tile_X65Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101010101010010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X66Y32, nonlinear_LMDPL
constant Tile_X66Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000101010100000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000011001100110011000000000000000000010001000100010";
--X67Y32, linear_LMDPL
constant Tile_X67Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000111111111010101011111111000000000000000010101010000000001010101010101010000000000000000000000000101010100000000000000000001000100010001000000000000000001010101010101010";
--X68Y32, linear_LMDPL
constant Tile_X68Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000011001100110011";
--X69Y32, nonlinear_LMDPL
constant Tile_X69Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101001010101000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y32, linear_LMDPL
constant Tile_X70Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001010101010101010";
--X71Y32, linear_LMDPL
constant Tile_X71Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000101010100000000000000000011101110111011110111011101110110000000000000000";
--X72Y32, nonlinear_LMDPL
constant Tile_X72Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X73Y32, linear_LMDPL
constant Tile_X73Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000010001000100010";
--X74Y32, linear_LMDPL
constant Tile_X74Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X75Y32, nonlinear_LMDPL
constant Tile_X75Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000100010001000100000000101010100010001000100010000000000000000000000000000000001100110011001100";
--X76Y32, linear_LMDPL
constant Tile_X76Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X77Y32, linear_LMDPL
constant Tile_X77Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000000000000000000";
--X78Y32, ctrl_to_sec
constant Tile_X78Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y32, combined_WDDL
constant Tile_X79Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011100000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110000000000000000000000000101010110100000101010100000101001000100000000001111111100000000";
--X80Y32, combined_WDDL
constant Tile_X80Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000011110000000000000000111100000000101000000000000000000000000000000101010100000000000010101010000011001100000000001011101100000000";
--X81Y32, ctrl_IO
constant Tile_X81Y32_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y33, W_IO_custom
constant Tile_X0Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y33, linear_LMDPL
constant Tile_X1Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000101010101010101011111111000000001111111100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X2Y33, linear_LMDPL
constant Tile_X2Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101100110011001100000000000000000";
--X3Y33, nonlinear_LMDPL
constant Tile_X3Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X4Y33, linear_LMDPL
constant Tile_X4Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000001010101010101010101010100000000000000000001000100010001000000000000000010011001100110010000000000000000";
--X5Y33, linear_LMDPL
constant Tile_X5Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000010011001100110010000000000000000";
--X6Y33, nonlinear_LMDPL
constant Tile_X6Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000";
--X7Y33, linear_LMDPL
constant Tile_X7Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000111111111010101000000000010101010101010100000000101010101001100110011001000000000000000000010001000100010000000000000000";
--X8Y33, linear_LMDPL
constant Tile_X8Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100000000010101010000000000000000000000000000000000101010111111111000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000000010001000100010000000000000000";
--X9Y33, nonlinear_LMDPL
constant Tile_X9Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000100010001000100100010001000100000000000000000";
--X10Y33, linear_LMDPL
constant Tile_X10Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000111111110101010101010101010101011010101000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001011101110111011";
--X11Y33, linear_LMDPL
constant Tile_X11Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000101010100000000000000000000000000101010101010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X12Y33, nonlinear_LMDPL
constant Tile_X12Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010111111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101010101010101010100000000000000001100110011001100000000000000000001000100010001000000000000000000";
--X13Y33, linear_LMDPL
constant Tile_X13Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X14Y33, linear_LMDPL
constant Tile_X14Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X15Y33, nonlinear_LMDPL
constant Tile_X15Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000001001100110011001";
--X16Y33, linear_LMDPL
constant Tile_X16Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X17Y33, linear_LMDPL
constant Tile_X17Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X18Y33, nonlinear_LMDPL
constant Tile_X18Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000011001100110011001000100010001000000000000000000";
--X19Y33, linear_LMDPL
constant Tile_X19Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000001010101000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X20Y33, linear_LMDPL
constant Tile_X20Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X21Y33, nonlinear_LMDPL
constant Tile_X21Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X22Y33, linear_LMDPL
constant Tile_X22Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X23Y33, linear_LMDPL
constant Tile_X23Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X24Y33, nonlinear_LMDPL
constant Tile_X24Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000011111111010001000100010000000000101010100000000000000000011101110111011110101010101010100000000000000000";
--X25Y33, linear_LMDPL
constant Tile_X25Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000001100110011001110101010101010100000000000000000";
--X26Y33, linear_LMDPL
constant Tile_X26Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000111111111001100110011001000000000000000010101010101010100000000000000000";
--X27Y33, nonlinear_LMDPL
constant Tile_X27Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000010101010010001000100010000000000000000000000000000000000110011001100110011001100110011000000000000000000";
--X28Y33, linear_LMDPL
constant Tile_X28Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000001101110111011101000000000000000000000000000000001100110011001100";
--X29Y33, linear_LMDPL
constant Tile_X29Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000100010001000100000000000000000000011001100110011";
--X30Y33, nonlinear_LMDPL
constant Tile_X30Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000010001000100010";
--X31Y33, linear_LMDPL
constant Tile_X31Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000100010001000111111111000000000101010101010101000000000000000000000000000000000000000000000000";
--X32Y33, linear_LMDPL
constant Tile_X32Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000110011001100110000000000000000001000100010001000";
--X33Y33, nonlinear_LMDPL
constant Tile_X33Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X34Y33, linear_LMDPL
constant Tile_X34Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X35Y33, linear_LMDPL
constant Tile_X35Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000010001000100010";
--X36Y33, nonlinear_LMDPL
constant Tile_X36Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000011001100110011";
--X37Y33, linear_LMDPL
constant Tile_X37Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000010101010000000000000000000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X38Y33, linear_LMDPL
constant Tile_X38Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000001100110011001101110111011101110000000000000000";
--X39Y33, nonlinear_LMDPL
constant Tile_X39Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y33, linear_LMDPL
constant Tile_X40Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010000000000000000010101010101010100000000000000001010101010101010000000000000000011011101110111010000000000000000";
--X41Y33, linear_LMDPL
constant Tile_X41Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101111111100000000000000001111111100000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X42Y33, nonlinear_LMDPL
constant Tile_X42Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101000000000101010101010101010101010000000000000000000000000000000000000000010101010000100010001000100000000000000000001000100010001000000000000000000000000000000000100010001000100";
--X43Y33, linear_LMDPL
constant Tile_X43Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010101010101010110101010101010100000000000000000";
--X44Y33, linear_LMDPL
constant Tile_X44Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010101010100000000011111111101010100000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X45Y33, nonlinear_LMDPL
constant Tile_X45Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000101010101010101000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X46Y33, linear_LMDPL
constant Tile_X46Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000001010101000000000000000000101010100000000010001000100010001010101000000000000000000000000111011101110111010101010101010100000000000000000";
--X47Y33, linear_LMDPL
constant Tile_X47Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000010101010101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001111111111111111";
--X48Y33, nonlinear_LMDPL
constant Tile_X48Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000000000000010101011010101001010101000000000000000000000000000000000000000000000000100010001000100000000000000000000001000100010001";
--X49Y33, linear_LMDPL
constant Tile_X49Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000001111111110101010111111110000000010101010000000000000000010101010101010100101010101010101000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X50Y33, linear_LMDPL
constant Tile_X50Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000100010001000100000000000000001010101010101010000000000000000000000000000000001100110011001100";
--X51Y33, nonlinear_LMDPL
constant Tile_X51Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101010101000000000101010100000000000000000000000000000000000000000111111111010101010101010000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000000000001100110011001100000000000000001001100110011001";
--X52Y33, linear_LMDPL
constant Tile_X52Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010101010100000000000000000101010100000000000000000000000000000000010101010000000001010101010101010000000000000000011111111000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000010001000100010";
--X53Y33, linear_LMDPL
constant Tile_X53Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010101011010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110110111011101110110000000000000000";
--X54Y33, nonlinear_LMDPL
constant Tile_X54Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000111111110000000000000000000000000000000010101010000000000101010100000000000000000000000000000000010101010000000000000000000100010001000100000000000000001000100010001000";
--X55Y33, linear_LMDPL
constant Tile_X55Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000011111111010101010000000000000000101010100000000000000000101010100000000001010101101010100101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X56Y33, linear_LMDPL
constant Tile_X56Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000010101011010101010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X57Y33, nonlinear_LMDPL
constant Tile_X57Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000110011001100110000000000000000001000100010001000000000000000000";
--X58Y33, linear_LMDPL
constant Tile_X58Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000010101010000000010101010000000000000000000000000010101010101010100000000101010100000000000000000010101011010101010101010010001000100010010101010010101010000000000000000110111011101110111011101110111010000000000000000";
--X59Y33, linear_LMDPL
constant Tile_X59Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000010101010000000000000000010101010000000000000000011111111101010101010101010101010010001000100010011111111010101010000000000000000010101010101010100000000000000000000000000000000";
--X60Y33, nonlinear_LMDPL
constant Tile_X60Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000011111111000000001010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001001100110011001";
--X61Y33, linear_LMDPL
constant Tile_X61Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000101010100000000000000000000000001010101101010101010101000000000010101010101010110101010101010100000000000000000000000000000000011111111111111110000000000000000";
--X62Y33, linear_LMDPL
constant Tile_X62Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000001010101101010100000000000000000111111110000000010101010101010100101010110101010000000000000000010101010000000000000000011111111000100010001000100000000101010100100010001000100000000000000000000000000000000001000100010001000";
--X63Y33, nonlinear_LMDPL
constant Tile_X63Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000000000101010100000000000000000000000010101010000000000000000000000000101010101010101001010101000100010001000100000000000000000110011001100110000000000000000000000000000000000101010101010101";
--X64Y33, linear_LMDPL
constant Tile_X64Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010101010101001010101010001000100010000000000101010100000000000000000100010001000100010001000100010000000000000000000";
--X65Y33, linear_LMDPL
constant Tile_X65Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000111111111010101010101010010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X66Y33, nonlinear_LMDPL
constant Tile_X66Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000101010101010101";
--X67Y33, linear_LMDPL
constant Tile_X67Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000111111111010101010101010000000000000000000000000000000001010101010101010000100010001000100000000101010101000100010001000000000000000000000000000000000001010101010101010";
--X68Y33, linear_LMDPL
constant Tile_X68Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000010101010101010100000000010101010010101010101010100000000101010101011101110111011000000000000000001010101010101010000000000000000";
--X69Y33, nonlinear_LMDPL
constant Tile_X69Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X70Y33, linear_LMDPL
constant Tile_X70Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X71Y33, linear_LMDPL
constant Tile_X71Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000101010101010101";
--X72Y33, nonlinear_LMDPL
constant Tile_X72Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X73Y33, linear_LMDPL
constant Tile_X73Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101011111111000000000000000000000000101010100000000000000000110011001100110000000000000000001011101110111011";
--X74Y33, linear_LMDPL
constant Tile_X74Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000001010101000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001000100010001000";
--X75Y33, nonlinear_LMDPL
constant Tile_X75Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010101010101000000000000100010001000100000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X76Y33, linear_LMDPL
constant Tile_X76Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010010001000100010000000000000000000000000000000000001000100010001010001000100010000000000000000000";
--X77Y33, linear_LMDPL
constant Tile_X77Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100110101010101010100000000000000000";
--X78Y33, ctrl_to_sec
constant Tile_X78Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000";
--X79Y33, combined_WDDL
constant Tile_X79Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000101010101111101011111111000000000100010000000000";
--X80Y33, combined_WDDL
constant Tile_X80Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000101000000000000010100000000000000000000000000101010100000000111100001010000010011001000000001100110000000000";
--X81Y33, ctrl_IO
constant Tile_X81Y33_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y34, W_IO_custom
constant Tile_X0Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y34, linear_LMDPL
constant Tile_X1Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000101010100000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X2Y34, linear_LMDPL
constant Tile_X2Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000001010101000000000101010111111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X3Y34, nonlinear_LMDPL
constant Tile_X3Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001";
--X4Y34, linear_LMDPL
constant Tile_X4Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X5Y34, linear_LMDPL
constant Tile_X5Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100101010100000000010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X6Y34, nonlinear_LMDPL
constant Tile_X6Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010000000000000000000000000000000010101010000000000101010100000000000000000000000001010101010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X7Y34, linear_LMDPL
constant Tile_X7Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000011111111101010100000000000000000010001000100010000000000000000000000000000000000001100110011001100100010001000100000000000000000";
--X8Y34, linear_LMDPL
constant Tile_X8Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010101010101010101010000000000101010100000000000000001111111110101010010001000100010000000000000000000000000000000000001100110011001110101010101010100000000000000000";
--X9Y34, nonlinear_LMDPL
constant Tile_X9Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000010111011101110110000000000000000";
--X10Y34, linear_LMDPL
constant Tile_X10Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101010101010101010101010101000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000001100110011001100";
--X11Y34, linear_LMDPL
constant Tile_X11Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010110101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000010001000100010";
--X12Y34, nonlinear_LMDPL
constant Tile_X12Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000001010101000000000101010100000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001100110011001100000000000000000000000000000000001001100110011001";
--X13Y34, linear_LMDPL
constant Tile_X13Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100110111011101110110000000000000000";
--X14Y34, linear_LMDPL
constant Tile_X14Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X15Y34, nonlinear_LMDPL
constant Tile_X15Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X16Y34, linear_LMDPL
constant Tile_X16Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X17Y34, linear_LMDPL
constant Tile_X17Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X18Y34, nonlinear_LMDPL
constant Tile_X18Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y34, linear_LMDPL
constant Tile_X19Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000110011001100110001010101010101010000000000000000";
--X20Y34, linear_LMDPL
constant Tile_X20Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000011111111000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X21Y34, nonlinear_LMDPL
constant Tile_X21Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010101010101101010100000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000011001100110011000000000000000000001000100010001";
--X22Y34, linear_LMDPL
constant Tile_X22Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101111111100000000010001000100010000000000000000000000000000000000010001000100010011111111111111110000000000000000";
--X23Y34, linear_LMDPL
constant Tile_X23Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000111111110000000000000000010001000100010010001000100010000000000000000000";
--X24Y34, nonlinear_LMDPL
constant Tile_X24Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111110101010010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X25Y34, linear_LMDPL
constant Tile_X25Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000000000000000000010101010101010100000000000000000";
--X26Y34, linear_LMDPL
constant Tile_X26Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000010101010000000001010101010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X27Y34, nonlinear_LMDPL
constant Tile_X27Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001100110011001100000000000000000000000000000000000101010101010101";
--X28Y34, linear_LMDPL
constant Tile_X28Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111010101010000000010101010000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000111011101110111";
--X29Y34, linear_LMDPL
constant Tile_X29Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X30Y34, nonlinear_LMDPL
constant Tile_X30Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X31Y34, linear_LMDPL
constant Tile_X31Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000001011101110111011";
--X32Y34, linear_LMDPL
constant Tile_X32Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X33Y34, nonlinear_LMDPL
constant Tile_X33Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y34, linear_LMDPL
constant Tile_X34Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000011001100110011";
--X35Y34, linear_LMDPL
constant Tile_X35Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X36Y34, nonlinear_LMDPL
constant Tile_X36Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000101010101010101";
--X37Y34, linear_LMDPL
constant Tile_X37Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010101111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X38Y34, linear_LMDPL
constant Tile_X38Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X39Y34, nonlinear_LMDPL
constant Tile_X39Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y34, linear_LMDPL
constant Tile_X40Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000101010100000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010101010101010111001100110011000000000000000000";
--X41Y34, linear_LMDPL
constant Tile_X41Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001100110011001100";
--X42Y34, nonlinear_LMDPL
constant Tile_X42Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100101010100000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X43Y34, linear_LMDPL
constant Tile_X43Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010110101010000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X44Y34, linear_LMDPL
constant Tile_X44Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100101010110101010000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000110011001100110011001100110011000000000000000000";
--X45Y34, nonlinear_LMDPL
constant Tile_X45Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000101010100101010100000000000000000000000000000000000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X46Y34, linear_LMDPL
constant Tile_X46Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000011111111000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X47Y34, linear_LMDPL
constant Tile_X47Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000100010001000100000000101010100100010001000100000000000000000000000000000000001011101110111011";
--X48Y34, nonlinear_LMDPL
constant Tile_X48Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000001111111100000000000000001010101010101010010101010101010100000000000000000001000100010001000000000000000011001100110011000000000000000000";
--X49Y34, linear_LMDPL
constant Tile_X49Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000001010101010101010101010100000000010101010000000000000000000000000101010100101010111111111010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X50Y34, linear_LMDPL
constant Tile_X50Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000000100010001000100100010001000100000000000000000";
--X51Y34, nonlinear_LMDPL
constant Tile_X51Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000000111111111010101000000000000000000101010110101010000000000000000010101010000000001010101000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000001000100010001";
--X52Y34, linear_LMDPL
constant Tile_X52Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101010101000000000000000000000000000000000";
--X53Y34, linear_LMDPL
constant Tile_X53Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000101010100101010110101010000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X54Y34, nonlinear_LMDPL
constant Tile_X54Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001100110011001100";
--X55Y34, linear_LMDPL
constant Tile_X55Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101101010100000000000000000101010100101010100000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000110011001100110000000000000000000101010101010101";
--X56Y34, linear_LMDPL
constant Tile_X56Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000101010100000000000000000000000010101010000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X57Y34, nonlinear_LMDPL
constant Tile_X57Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010101010101010101010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X58Y34, linear_LMDPL
constant Tile_X58Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000111111110000000000000000000000001010101011111111000000000000000000000000000000001010101010101010000100010001000100000000000000001010101010101010000000000000000000000000000000001101110111011101";
--X59Y34, linear_LMDPL
constant Tile_X59Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010100101010100000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000101010110101010000000000000000011111111000000001010101010101010010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X60Y34, nonlinear_LMDPL
constant Tile_X60Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101000000000101010101010101010101010000000000000000000000000000000001010101000000000010101010101010100000000101010101110111011101110000000000000000000000000000000000000000000000000";
--X61Y34, linear_LMDPL
constant Tile_X61Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X62Y34, linear_LMDPL
constant Tile_X62Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101011010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010101010101001010101000000000000000000000000000000000000000010101010010101010101010100000000101010101010101010101010000000000000000001000100010001000000000000000000";
--X63Y34, nonlinear_LMDPL
constant Tile_X63Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010101010101010101010000100010001000100000000101010101001100110011001000000000000000000000000000000000011001100110011";
--X64Y34, linear_LMDPL
constant Tile_X64Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010101111111100000000000000001010101000000000101010101010101000000000000000000000000010101010101010101010101001010101000100010001000111111111000000001010101010101010000000000000000000000000000000001000100010001000";
--X65Y34, linear_LMDPL
constant Tile_X65Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000010101010111111110000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010101010101010101010010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X66Y34, nonlinear_LMDPL
constant Tile_X66Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000010101010000100010001000100000000101010101011101110111011000000000000000000000000000000000000000000000000";
--X67Y34, linear_LMDPL
constant Tile_X67Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000101010100101010111111111000000000000000010101010101010101010101011111111000000000000000011111111101010100000000000000000000000000000000000000000000000001000100010001000";
--X68Y34, linear_LMDPL
constant Tile_X68Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000010101010000000000000000010101010000000000000000000000000001000100010001000000000000000000100010001000100";
--X69Y34, nonlinear_LMDPL
constant Tile_X69Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010110101010000000000000000010101010000000001010101000000000000100010001000100000000010101010000000000000000000000000000000000000000000000001000100010001000";
--X70Y34, linear_LMDPL
constant Tile_X70Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X71Y34, linear_LMDPL
constant Tile_X71Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X72Y34, nonlinear_LMDPL
constant Tile_X72Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101111111100000000010101010101010100000000000000000100010001000100000000000000000001010101010101010000000000000000";
--X73Y34, linear_LMDPL
constant Tile_X73Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000010101010000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X74Y34, linear_LMDPL
constant Tile_X74Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X75Y34, nonlinear_LMDPL
constant Tile_X75Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000101010101111111100000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X76Y34, linear_LMDPL
constant Tile_X76Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000011111111000000000000000010101010010101010000000010101010010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X77Y34, linear_LMDPL
constant Tile_X77Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X78Y34, ctrl_to_sec
constant Tile_X78Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000";
--X79Y34, combined_WDDL
constant Tile_X79Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100001111101010101010101011001100000000000000000000000000";
--X80Y34, combined_WDDL
constant Tile_X80Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000000101000000000000000000000000000000000000000000000111100000000101000000000000000000000000000000101010100000000000000001010000011011101000000001011101100000000";
--X81Y34, ctrl_IO
constant Tile_X81Y34_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y35, W_IO_custom
constant Tile_X0Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y35, linear_LMDPL
constant Tile_X1Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101000000000000000001010101000000000101010100000000001010101000000000000000010101010010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X2Y35, linear_LMDPL
constant Tile_X2Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101010101010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110010011001100110010000000000000000";
--X3Y35, nonlinear_LMDPL
constant Tile_X3Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000010101010000000010101010010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X4Y35, linear_LMDPL
constant Tile_X4Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111110101010000000001010101000000000101010100000000010101010000000000000000000000000010101010000000000000000001000100010001000000000000000000011001100110011";
--X5Y35, linear_LMDPL
constant Tile_X5Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010101010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X6Y35, nonlinear_LMDPL
constant Tile_X6Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X7Y35, linear_LMDPL
constant Tile_X7Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000001010101010101010101010100000000101010101011101110111011000000000000000010011001100110010000000000000000";
--X8Y35, linear_LMDPL
constant Tile_X8Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101011111111110101010010101010000000000000000000000000000000001010101101010100000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000010011001100110010000000000000000";
--X9Y35, nonlinear_LMDPL
constant Tile_X9Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X10Y35, linear_LMDPL
constant Tile_X10Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000101010110101010101010101111111100000000000000001010101000000000000000000000000010101010010101010101010100000000000000001001100110011001000000000000000011001100110011000000000000000000";
--X11Y35, linear_LMDPL
constant Tile_X11Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X12Y35, nonlinear_LMDPL
constant Tile_X12Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100";
--X13Y35, linear_LMDPL
constant Tile_X13Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000111111110000000010101010000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X14Y35, linear_LMDPL
constant Tile_X14Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111110101010000000000000000000000000000000001111111100000000000000000000000010101010010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X15Y35, nonlinear_LMDPL
constant Tile_X15Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X16Y35, linear_LMDPL
constant Tile_X16Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000010001000100010000000000000000000000000000000000100110011001100100100010001000100000000000000000";
--X17Y35, linear_LMDPL
constant Tile_X17Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001011101110111011";
--X18Y35, nonlinear_LMDPL
constant Tile_X18Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000001000100010001";
--X19Y35, linear_LMDPL
constant Tile_X19Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X20Y35, linear_LMDPL
constant Tile_X20Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X21Y35, nonlinear_LMDPL
constant Tile_X21Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000111111111010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001101110111011101";
--X22Y35, linear_LMDPL
constant Tile_X22Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101001010101000000000101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X23Y35, linear_LMDPL
constant Tile_X23Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X24Y35, nonlinear_LMDPL
constant Tile_X24Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010101111111110101010000000000000000000000000101010100000000000000000011001100110011000000000000000000100010001000100";
--X25Y35, linear_LMDPL
constant Tile_X25Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X26Y35, linear_LMDPL
constant Tile_X26Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000011111111101010100000000000000000000100010001000111111111101010100010001000100010000000000000000000000000000000000110011001100110";
--X27Y35, nonlinear_LMDPL
constant Tile_X27Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000101010101010101010101010000000000000000000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000010011001100110010000000000000000";
--X28Y35, linear_LMDPL
constant Tile_X28Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001101110111011101";
--X29Y35, linear_LMDPL
constant Tile_X29Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000011111111000000000000000010101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X30Y35, nonlinear_LMDPL
constant Tile_X30Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011";
--X31Y35, linear_LMDPL
constant Tile_X31Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000010101010000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X32Y35, linear_LMDPL
constant Tile_X32Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000111111111111111110101010101010100000000000000000";
--X33Y35, nonlinear_LMDPL
constant Tile_X33Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X34Y35, linear_LMDPL
constant Tile_X34Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X35Y35, linear_LMDPL
constant Tile_X35Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X36Y35, nonlinear_LMDPL
constant Tile_X36Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000010001000100010";
--X37Y35, linear_LMDPL
constant Tile_X37Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X38Y35, linear_LMDPL
constant Tile_X38Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X39Y35, nonlinear_LMDPL
constant Tile_X39Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X40Y35, linear_LMDPL
constant Tile_X40Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000110111011101110100000000000000000101010101010101";
--X41Y35, linear_LMDPL
constant Tile_X41Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111110101010101010100101010111111111010101010000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X42Y35, nonlinear_LMDPL
constant Tile_X42Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000010011001100110010000000000000000";
--X43Y35, linear_LMDPL
constant Tile_X43Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010100000000000000000010101010101010100000000010101010100010001000100000000000000000011001100110011000000000000000000";
--X44Y35, linear_LMDPL
constant Tile_X44Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101001010101101010100101010100000000000000000101010100000000101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000011011101110111010000000000000000";
--X45Y35, nonlinear_LMDPL
constant Tile_X45Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000101010100101010100000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000011101110111011100000000000000001000100010001000";
--X46Y35, linear_LMDPL
constant Tile_X46Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000001111111100000000000000001010101000000000010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X47Y35, linear_LMDPL
constant Tile_X47Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X48Y35, nonlinear_LMDPL
constant Tile_X48Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000100010001000100001110111011101110000000000000000";
--X49Y35, linear_LMDPL
constant Tile_X49Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001010101000000000101010100101010110101010000000000000000010101010101010100101010111111111010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X50Y35, linear_LMDPL
constant Tile_X50Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010101010101000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000100010001000100";
--X51Y35, nonlinear_LMDPL
constant Tile_X51Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100101010110101010101010101111111100000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000000010001000100010";
--X52Y35, linear_LMDPL
constant Tile_X52Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010000000000000000000000101010100101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101111111110101010100000000000000000000000010101010010101010000000000000000010001000100010000000000000000000000000000000000111011101110111000000000000000000000000000000000";
--X53Y35, linear_LMDPL
constant Tile_X53Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000111111111010101010101010000000000000000000000000000000000101010110101010010001000100010000000000010101010000000000000000000000000000000010111011101110110000000000000000";
--X54Y35, nonlinear_LMDPL
constant Tile_X54Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010101010101001010101000000000000000010101010000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011";
--X55Y35, linear_LMDPL
constant Tile_X55Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X56Y35, linear_LMDPL
constant Tile_X56Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000111111111010101010101010000000000000000011111111101010100000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X57Y35, nonlinear_LMDPL
constant Tile_X57Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010111111111010101010101010000000000000000001010101000000001010101001010101000000000000000000000000101010100000000000000000110011001100110000000000000000001010101010101010";
--X58Y35, linear_LMDPL
constant Tile_X58Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000010101010010101010000000000000000000000001010101000000000000000000000000011111111000000001010101000000000000100010001000100000000010101011000100010001000000000000000000000000000000000001011101110111011";
--X59Y35, linear_LMDPL
constant Tile_X59Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000101010100000000000000000000000011111111000000001010101010101010010101010101010100000000101010101000100010001000000000000000000011011101110111010000000000000000";
--X60Y35, nonlinear_LMDPL
constant Tile_X60Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000101010101010101000000000000000001111111101010101000000000000000001010101111111110000000010101010000000001010101000000000101010100101010110101010000000000000000000000000010101011010101001010101010101010101010100000000000000001101110111011101000000000000000001110111011101110000000000000000";
--X61Y35, linear_LMDPL
constant Tile_X61Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X62Y35, linear_LMDPL
constant Tile_X62Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010111111110101010110101010000000000000000010101010000000000000000010101010000100010001000100000000101010101101110111011101000000000000000000000000000000001000100010001000";
--X63Y35, nonlinear_LMDPL
constant Tile_X63Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000101010100000000000000000000100010001000110101010101010100000000000000000";
--X64Y35, linear_LMDPL
constant Tile_X64Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000101010100101010100000000000000000000000000000000101010101010101001010101000100010001000100000000101010100111011101110111000000000000000000000000000000000101010101010101";
--X65Y35, linear_LMDPL
constant Tile_X65Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101001010101111111110000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000001010101000100010001000100000000010101011100110011001100000000000000000000000000000000001000100010001000";
--X66Y35, nonlinear_LMDPL
constant Tile_X66Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000101010101010101";
--X67Y35, linear_LMDPL
constant Tile_X67Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111111111110101010000000001010101000000000010101011010101010101010000000000000000000000000101010101010101000000000000100010001000100000000010101011010101010101010000000000000000000000000000000001000100010001000";
--X68Y35, linear_LMDPL
constant Tile_X68Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000010101010010101010101010100000000000000001101110111011101000000000000000000100010001000100000000000000000";
--X69Y35, nonlinear_LMDPL
constant Tile_X69Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000010101010111111110000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X70Y35, linear_LMDPL
constant Tile_X70Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000101010101010101";
--X71Y35, linear_LMDPL
constant Tile_X71Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000010001000100010010101010101010100000000000000000";
--X72Y35, nonlinear_LMDPL
constant Tile_X72Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111101010100000000000000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X73Y35, linear_LMDPL
constant Tile_X73Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X74Y35, linear_LMDPL
constant Tile_X74Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000101010100000000000000000000100010001000100110011001100110000000000000000";
--X75Y35, nonlinear_LMDPL
constant Tile_X75Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101011111111010101010101010100000000101010100101010101010101000000000000000010001000100010000000000000000000";
--X76Y35, linear_LMDPL
constant Tile_X76Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010101010101010101010000100010001000100000000010101011000100010001000000000000000000000000000000000000011001100110011";
--X77Y35, linear_LMDPL
constant Tile_X77Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X78Y35, ctrl_to_sec
constant Tile_X78Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000001011111000000000000000000000000000000000000000000001111000000000000000000000000";
--X79Y35, combined_WDDL
constant Tile_X79Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001111000000000000101010100000000000000000000000000101010100001010101010100000101010111011000000000011001100000000";
--X80Y35, combined_WDDL
constant Tile_X80Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000101010100000000000011110000000010111011000000001001100100000000";
--X81Y35, ctrl_IO
constant Tile_X81Y35_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y36, W_IO_custom
constant Tile_X0Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y36, linear_LMDPL
constant Tile_X1Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000001010101001010101000000000000000000000000010101010000000010101010010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X2Y36, linear_LMDPL
constant Tile_X2Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110000110011001100110000000000000000";
--X3Y36, nonlinear_LMDPL
constant Tile_X3Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X4Y36, linear_LMDPL
constant Tile_X4Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000111111111010101000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X5Y36, linear_LMDPL
constant Tile_X5Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001000100010001000000000000000000000110011001100110000000000000000";
--X6Y36, nonlinear_LMDPL
constant Tile_X6Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000010101010010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X7Y36, linear_LMDPL
constant Tile_X7Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000010101010010101010101010100000000000000000111011101110111000000000000000011001100110011000000000000000000";
--X8Y36, linear_LMDPL
constant Tile_X8Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010111111111000000000000000000000000000000000000000010101010010101010000000010101010000000000000000000000000111111111010101000000000010101010101010100000000000000000110011001100110000000000000000010001000100010000000000000000000";
--X9Y36, nonlinear_LMDPL
constant Tile_X9Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000001000100010001000000000000000000110011001100110000000000000000";
--X10Y36, linear_LMDPL
constant Tile_X10Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010000000001111111111111111000000000000000010101010101010100000000000000000000000000101010100000000111111110000000000000000010101010101010100000000000000000101010101010101000000000000000010101010101010100000000000000000";
--X11Y36, linear_LMDPL
constant Tile_X11Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X12Y36, nonlinear_LMDPL
constant Tile_X12Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101100110011001100110000000000000000";
--X13Y36, linear_LMDPL
constant Tile_X13Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X14Y36, linear_LMDPL
constant Tile_X14Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000101110111011101100000000000000001110111011101110";
--X15Y36, nonlinear_LMDPL
constant Tile_X15Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X16Y36, linear_LMDPL
constant Tile_X16Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100110111011101110110000000000000000";
--X17Y36, linear_LMDPL
constant Tile_X17Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X18Y36, nonlinear_LMDPL
constant Tile_X18Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000011001100110011000100010001000100000000000000000";
--X19Y36, linear_LMDPL
constant Tile_X19Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000001000100010001000000000000000000000000000000000";
--X20Y36, linear_LMDPL
constant Tile_X20Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000011111111010101010101010100000000000000001101110111011101000000000000000001110111011101110000000000000000";
--X21Y36, nonlinear_LMDPL
constant Tile_X21Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111010101010000000001010101000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000100010001000100010011001100110010000000000000000";
--X22Y36, linear_LMDPL
constant Tile_X22Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000001111111100000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010001000100010011111111000000000000000000000000111111111111111100100010001000100000000000000000";
--X23Y36, linear_LMDPL
constant Tile_X23Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000101010101110111011101110000000000000000000000000000000000011001100110011";
--X24Y36, nonlinear_LMDPL
constant Tile_X24Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101010101010000100010001000100000000000000001001100110011001000000000000000000000000000000001010101010101010";
--X25Y36, linear_LMDPL
constant Tile_X25Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000010101010101010101000100010001000000000000000000";
--X26Y36, linear_LMDPL
constant Tile_X26Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X27Y36, nonlinear_LMDPL
constant Tile_X27Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101011111111000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110010001000100010000000000000000000";
--X28Y36, linear_LMDPL
constant Tile_X28Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X29Y36, linear_LMDPL
constant Tile_X29Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000100010001000100000000000000000001100110011001100";
--X30Y36, nonlinear_LMDPL
constant Tile_X30Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000001010101000000000010001000100010000000000000000000000000000000000100010001000100011011101110111010000000000000000";
--X31Y36, linear_LMDPL
constant Tile_X31Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000000000000000000010101010010101010101010110101010000000000101010101010101000000000000000011111111111111110000000000000000";
--X32Y36, linear_LMDPL
constant Tile_X32Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X33Y36, nonlinear_LMDPL
constant Tile_X33Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X34Y36, linear_LMDPL
constant Tile_X34Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X35Y36, linear_LMDPL
constant Tile_X35Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X36Y36, nonlinear_LMDPL
constant Tile_X36Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000101010101010101";
--X37Y36, linear_LMDPL
constant Tile_X37Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010111111111000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X38Y36, linear_LMDPL
constant Tile_X38Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X39Y36, nonlinear_LMDPL
constant Tile_X39Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X40Y36, linear_LMDPL
constant Tile_X40Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001110111011101110000000000000000";
--X41Y36, linear_LMDPL
constant Tile_X41Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000010101010101010101010101010101010000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X42Y36, nonlinear_LMDPL
constant Tile_X42Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X43Y36, linear_LMDPL
constant Tile_X43Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000011111111000000000000000000000000010001000100010011111111000000000000000000000000010001000100010001010101010101010000000000000000";
--X44Y36, linear_LMDPL
constant Tile_X44Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000000100010001000100";
--X45Y36, nonlinear_LMDPL
constant Tile_X45Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000111111110000000000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000101010100000000010001000100010000000000010101010000000000000000000100010001000101010101010101010000000000000000";
--X46Y36, linear_LMDPL
constant Tile_X46Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010101010101000000000000000000000000010101010000000000000000010101010000000001010101000000000010001000100010001010101000000000000000000000000011001100110011001000100010001000000000000000000";
--X47Y36, linear_LMDPL
constant Tile_X47Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000001010101010101010000000000000000000000000000000000000000000000000101010100000000111111110000000000000000010101010101010100000000000100010001000100000000101010100101010101010101000000000000000000000000000000001000100010001000";
--X48Y36, nonlinear_LMDPL
constant Tile_X48Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000111111110000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000101010110101010010101010101010100000000000000000000000000000000000000000000000000010001000100010000000000000000";
--X49Y36, linear_LMDPL
constant Tile_X49Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101000000000101010101010101001010101000000000000000000000000000000000101010110101010010001000100010000000000000000000000000000000000101110111011101110101010101010100000000000000000";
--X50Y36, linear_LMDPL
constant Tile_X50Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010111111111000000000000000001010101101010101010101010101010010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X51Y36, nonlinear_LMDPL
constant Tile_X51Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000001010101111111110000000000000000000000001010101000000000010101010101010110101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X52Y36, linear_LMDPL
constant Tile_X52Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010110101010000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X53Y36, linear_LMDPL
constant Tile_X53Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101101010100000000000000000101010100000000000000000000000000000000001010101000000001010101010101010000000000000000000000000010101011010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X54Y36, nonlinear_LMDPL
constant Tile_X54Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000001010101101010101010101010101010000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X55Y36, linear_LMDPL
constant Tile_X55Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010110101010010101010000000000000000101010101010101000000000000000000101010100000000101010100000000000000000111111111010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X56Y36, linear_LMDPL
constant Tile_X56Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000000000000000000001010101010101010000000000101010110101010010101010000000010101010010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X57Y36, nonlinear_LMDPL
constant Tile_X57Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111101010101101010101010101010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X58Y36, linear_LMDPL
constant Tile_X58Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000010101010000000011111111000000001111111100000000101010100000000010101010000000001010101001010101101010100000000000000000101010100101010100000000010101010101010110101010000000000101010101010101000000000000000000100010001000100000000000000000";
--X59Y36, linear_LMDPL
constant Tile_X59Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010101010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000010101010010101010000000001010101000100010001000110101010000000001010101010101010000000000000000000000000000000001010101010101010";
--X60Y36, nonlinear_LMDPL
constant Tile_X60Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101010101010000000000000000000000000101010101010101010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000001000100010001";
--X61Y36, linear_LMDPL
constant Tile_X61Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000110101010000000000100010001000100000000000000000000000000000000000000000000000000";
--X62Y36, linear_LMDPL
constant Tile_X62Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000101010100000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000011111111111111110000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000001100110011001100";
--X63Y36, nonlinear_LMDPL
constant Tile_X63Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000001010101001010101000000000000000000000000101010100000000000000000111011101110111000000000000000000101010101010101";
--X64Y36, linear_LMDPL
constant Tile_X64Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000111111111010101010101010000000000000000010101010101010101010101000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X65Y36, linear_LMDPL
constant Tile_X65Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000001000100010001";
--X66Y36, nonlinear_LMDPL
constant Tile_X66Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000010101010101010100000000010101010011001100110011000000000000000001000100010001000000000000000000";
--X67Y36, linear_LMDPL
constant Tile_X67Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000011111111101010100000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000010101010101010100101010100000000010001000100010000000000101010100000000000000000011101110111011110001000100010000000000000000000";
--X68Y36, linear_LMDPL
constant Tile_X68Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X69Y36, nonlinear_LMDPL
constant Tile_X69Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000101010110101010000000000000000000000000101010100000000000000000110011001100110000000000000000000100010001000100";
--X70Y36, linear_LMDPL
constant Tile_X70Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000101010101010101";
--X71Y36, linear_LMDPL
constant Tile_X71Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000010101010010001000100010000000000101010100000000000000000111011101110111001000100010001000000000000000000";
--X72Y36, nonlinear_LMDPL
constant Tile_X72Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101101010100000000010101010010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X73Y36, linear_LMDPL
constant Tile_X73Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000011001100110011";
--X74Y36, linear_LMDPL
constant Tile_X74Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010101010101010100000000000000000101010101010101000000000000000000100010001000100000000000000000";
--X75Y36, nonlinear_LMDPL
constant Tile_X75Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010101111111100000000010101010101010100000000101010100000000000000000000000000000000001010101010101010000000000000000";
--X76Y36, linear_LMDPL
constant Tile_X76Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000001101110111011101000000000000000000000000000000000011001100110011";
--X77Y36, linear_LMDPL
constant Tile_X77Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000101010101101110111011101000000000000000010001000100010000000000000000000";
--X78Y36, ctrl_to_sec
constant Tile_X78Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000";
--X79Y36, combined_WDDL
constant Tile_X79Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000101000000000000000000000101000000000101010100000000000000000000000000101010100000000101000000000111111101110000000000100010000000000";
--X80Y36, combined_WDDL
constant Tile_X80Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y36, ctrl_IO
constant Tile_X81Y36_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y37, W_IO_custom
constant Tile_X0Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y37, linear_LMDPL
constant Tile_X1Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101011010101000000000000000001010101000000000101010100000000000000000000000001111111110101010010101010101010100000000000000001000100010001000000000000000000000010001000100010000000000000000";
--X2Y37, linear_LMDPL
constant Tile_X2Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X3Y37, nonlinear_LMDPL
constant Tile_X3Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111110101010000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X4Y37, linear_LMDPL
constant Tile_X4Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101101010100000000000000000000000000000000000000000000000001010101010101010000000001010101000000000101010100000000000000000010101010101010100000000101010100000000000000000000000000000000001000100010001000000000000000000";
--X5Y37, linear_LMDPL
constant Tile_X5Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000001010101000000000000000000000000000000000111111110000000000000000010101010101010100000000010101010000000000000000000000000000000010111011101110110000000000000000";
--X6Y37, nonlinear_LMDPL
constant Tile_X6Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010110101010010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X7Y37, linear_LMDPL
constant Tile_X7Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X8Y37, linear_LMDPL
constant Tile_X8Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X9Y37, nonlinear_LMDPL
constant Tile_X9Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X10Y37, linear_LMDPL
constant Tile_X10Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000010101010101010100000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000100010001000100000000000000000001100110011001100";
--X11Y37, linear_LMDPL
constant Tile_X11Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000010101010000000000101010100000000111111110000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000000010001000100010000000000000000";
--X12Y37, nonlinear_LMDPL
constant Tile_X12Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X13Y37, linear_LMDPL
constant Tile_X13Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000010101010000000010101010010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111";
--X14Y37, linear_LMDPL
constant Tile_X14Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X15Y37, nonlinear_LMDPL
constant Tile_X15Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000100010001000100000000010101010110011001100110000000000000000000000000000000000010001000100010";
--X16Y37, linear_LMDPL
constant Tile_X16Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000111011101110111010000000000000000";
--X17Y37, linear_LMDPL
constant Tile_X17Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X18Y37, nonlinear_LMDPL
constant Tile_X18Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X19Y37, linear_LMDPL
constant Tile_X19Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001000100010001000";
--X20Y37, linear_LMDPL
constant Tile_X20Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111111111100000000000000000101010101010101";
--X21Y37, nonlinear_LMDPL
constant Tile_X21Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111111010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X22Y37, linear_LMDPL
constant Tile_X22Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000011111111010101010101010101010101010101011010101010101010000000000000000010001000100010000000000000000000";
--X23Y37, linear_LMDPL
constant Tile_X23Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X24Y37, nonlinear_LMDPL
constant Tile_X24Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000110011001100110010001000100010000000000000000000";
--X25Y37, linear_LMDPL
constant Tile_X25Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000001111111100000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X26Y37, linear_LMDPL
constant Tile_X26Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000011111111000000000000000010101010010101010101010100000000000000001110111011101110000000000000000011011101110111010000000000000000";
--X27Y37, nonlinear_LMDPL
constant Tile_X27Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000001011101110111011";
--X28Y37, linear_LMDPL
constant Tile_X28Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X29Y37, linear_LMDPL
constant Tile_X29Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101001010101000000000000000010101010000000000101010110101010000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X30Y37, nonlinear_LMDPL
constant Tile_X30Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111101010100000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000001000100010001";
--X31Y37, linear_LMDPL
constant Tile_X31Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111101010101010101010101010000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000100010001000100010101010101010100000000000000000";
--X32Y37, linear_LMDPL
constant Tile_X32Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X33Y37, nonlinear_LMDPL
constant Tile_X33Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X34Y37, linear_LMDPL
constant Tile_X34Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X35Y37, linear_LMDPL
constant Tile_X35Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000011011101110111010000000000000000";
--X36Y37, nonlinear_LMDPL
constant Tile_X36Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000111011101110111000000000000000000100010001000100";
--X37Y37, linear_LMDPL
constant Tile_X37Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X38Y37, linear_LMDPL
constant Tile_X38Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X39Y37, nonlinear_LMDPL
constant Tile_X39Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y37, linear_LMDPL
constant Tile_X40Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000010101011111111110101010000000001010101000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X41Y37, linear_LMDPL
constant Tile_X41Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010110101010101010101010101000000000000000001010101011111111101010100000000000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X42Y37, nonlinear_LMDPL
constant Tile_X42Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X43Y37, linear_LMDPL
constant Tile_X43Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101010101010000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000010101010000000011111111000000000000000000000000101010100101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000000010001000100010";
--X44Y37, linear_LMDPL
constant Tile_X44Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000101010100000000101010101010101000000000000000000000000001010101000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X45Y37, nonlinear_LMDPL
constant Tile_X45Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100101010100000000000000000000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111000100010001000100000000000000000";
--X46Y37, linear_LMDPL
constant Tile_X46Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000001111111100000000010101010000000000000000101010101010101000000000000000000101010110101010000000000000000000000000000000000101010101010101010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X47Y37, linear_LMDPL
constant Tile_X47Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000010101010000000000000000110011001100110001000100010001000000000000000000";
--X48Y37, nonlinear_LMDPL
constant Tile_X48Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000101010100000000000000000000000000000000000000000010101011111111110101010101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110";
--X49Y37, linear_LMDPL
constant Tile_X49Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000001010101011111111101010101010101010101010000000000000000010101010000000000000000010101010010101010101010100000000010101010000000000000000000000000000000010111011101110110000000000000000";
--X50Y37, linear_LMDPL
constant Tile_X50Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101011111111000000000000000010101010101010101010101010101010010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X51Y37, nonlinear_LMDPL
constant Tile_X51Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000101010100000000000000000101010110101010000000000000000000000000000000000000000000000000010101010101010100000000101010101001100110011001000000000000000010101010101010100000000000000000";
--X52Y37, linear_LMDPL
constant Tile_X52Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000001111111100000000101010101010101010101010000100010001000100000000000000000011001100110011000000000000000000000000000000001000100010001000";
--X53Y37, linear_LMDPL
constant Tile_X53Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000101010101010101000000000000000000000000011111111101010101010101010101010010101010101010111111111010101011000100010001000000000000000000000000000000000000000000000000000";
--X54Y37, nonlinear_LMDPL
constant Tile_X54Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101111111111010101010101010000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000110011001100110000000000000000001111111111111111";
--X55Y37, linear_LMDPL
constant Tile_X55Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X56Y37, linear_LMDPL
constant Tile_X56Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000111111110000000000000000000000001010101000000000000000000101010110101010000000000000000010101010101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000101010110101010010001000100010000000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X57Y37, nonlinear_LMDPL
constant Tile_X57Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010000000000000000010101010010101010000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001000100010001000";
--X58Y37, linear_LMDPL
constant Tile_X58Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000101010110101010101010100000000000000000000000000000000011111111010101010101010100000000101010101101110111011101000000000000000011001100110011000000000000000000";
--X59Y37, linear_LMDPL
constant Tile_X59Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000101010100000000000000000000000010101010000000001010101000000000010101010000000000000000000000000101010100000000010101011010101000000000000000000000000010101010010101011010101000000000000100010001000100000000101010100000000000000000000000000000000000000000000000001101110111011101";
--X60Y37, nonlinear_LMDPL
constant Tile_X60Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000101010101010101000000000000000000000000000000001010101010101010000100010001000100000000010101010011001100110011000000000000000000000000000000000000000000000000";
--X61Y37, linear_LMDPL
constant Tile_X61Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000101010100000000000000000000100010001000100000000000000001100110011001100";
--X62Y37, linear_LMDPL
constant Tile_X62Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000001010101000000001111111110101010010101010000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010101100110011001100000000000000000001000100010001000000000000000000";
--X63Y37, nonlinear_LMDPL
constant Tile_X63Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000100110011001100100000000000000000000000000000000";
--X64Y37, linear_LMDPL
constant Tile_X64Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000101010110101010000000000000000000000000101010101010101000000000000100010001000100000000101010101111111111111111000000000000000000000000000000001010101010101010";
--X65Y37, linear_LMDPL
constant Tile_X65Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X66Y37, nonlinear_LMDPL
constant Tile_X66Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000001000100010001000";
--X67Y37, linear_LMDPL
constant Tile_X67Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010101010101000000000000000001010101000000000000000000101010111111111000000000000000000000000101010101010101000000000010001000100010000000000101010100000000000000000000000000000000000100010001000100000000000000000";
--X68Y37, linear_LMDPL
constant Tile_X68Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000101010101010101010101010010001000100010010101010000000000000000000000000000000000000000010001000100010000000000000000000";
--X69Y37, nonlinear_LMDPL
constant Tile_X69Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y37, linear_LMDPL
constant Tile_X70Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000000011001100110011000000000000000011011101110111010000000000000000";
--X71Y37, linear_LMDPL
constant Tile_X71Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000001010101011111111000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X72Y37, nonlinear_LMDPL
constant Tile_X72Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X73Y37, linear_LMDPL
constant Tile_X73Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X74Y37, linear_LMDPL
constant Tile_X74Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101011111111100000000000100010001000100000000101010101000100010001000000000000000000000000000000000000011001100110011";
--X75Y37, nonlinear_LMDPL
constant Tile_X75Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111101010100000000001010101000000000000000001010101101010100000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100";
--X76Y37, linear_LMDPL
constant Tile_X76Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100000000010101010000100010001000100000000101010101101110111011101000000000000000000000000000000000011001100110011";
--X77Y37, linear_LMDPL
constant Tile_X77Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101001010101010101010101010111111111010101010101010101010101000000000000000010101010101010100000000000000000";
--X78Y37, ctrl_to_sec
constant Tile_X78Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y37, combined_WDDL
constant Tile_X79Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000101000000000000000000000000000000000000000000000";
--X80Y37, combined_WDDL
constant Tile_X80Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000";
--X81Y37, ctrl_IO
constant Tile_X81Y37_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y38, W_IO_custom
constant Tile_X0Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y38, linear_LMDPL
constant Tile_X1Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000101010100000000000000000000000001111111110101010010101010101010100000000000000000101010101010101000000000000000010111011101110110000000000000000";
--X2Y38, linear_LMDPL
constant Tile_X2Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001011101110111011";
--X3Y38, nonlinear_LMDPL
constant Tile_X3Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000010101010010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X4Y38, linear_LMDPL
constant Tile_X4Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000100010001000100000000000000001001100110011001000000000000000000000000000000000001000100010001";
--X5Y38, linear_LMDPL
constant Tile_X5Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000000000001001100110011001000000000000000001000100010001000000000000000000";
--X6Y38, nonlinear_LMDPL
constant Tile_X6Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X7Y38, linear_LMDPL
constant Tile_X7Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X8Y38, linear_LMDPL
constant Tile_X8Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X9Y38, nonlinear_LMDPL
constant Tile_X9Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000010101010010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X10Y38, linear_LMDPL
constant Tile_X10Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111111010101001010101010101010000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001001100110011001";
--X11Y38, linear_LMDPL
constant Tile_X11Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001110011001100110010000000000000000";
--X12Y38, nonlinear_LMDPL
constant Tile_X12Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X13Y38, linear_LMDPL
constant Tile_X13Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001101110111011101";
--X14Y38, linear_LMDPL
constant Tile_X14Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000010101010101010100000000001010101000000001111111100000000000000000000000010101010010101010101010100000000000000000111011101110111000000000000000011101110111011100000000000000000";
--X15Y38, nonlinear_LMDPL
constant Tile_X15Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X16Y38, linear_LMDPL
constant Tile_X16Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X17Y38, linear_LMDPL
constant Tile_X17Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X18Y38, nonlinear_LMDPL
constant Tile_X18Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000100010001000100000000000000000";
--X19Y38, linear_LMDPL
constant Tile_X19Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X20Y38, linear_LMDPL
constant Tile_X20Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X21Y38, nonlinear_LMDPL
constant Tile_X21Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000010101010101010111111111000000001010101000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000001010101010101010";
--X22Y38, linear_LMDPL
constant Tile_X22Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X23Y38, linear_LMDPL
constant Tile_X23Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000100010001000100";
--X24Y38, nonlinear_LMDPL
constant Tile_X24Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001001100110011001";
--X25Y38, linear_LMDPL
constant Tile_X25Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000011111111000000001010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000011001100110011";
--X26Y38, linear_LMDPL
constant Tile_X26Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000011111111000000000000000011111111010101010101010100000000000000001010101010101010000000000000000011111111111111110000000000000000";
--X27Y38, nonlinear_LMDPL
constant Tile_X27Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000000100010001000100";
--X28Y38, linear_LMDPL
constant Tile_X28Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001100110011001100";
--X29Y38, linear_LMDPL
constant Tile_X29Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110101010110101010000000000000000001010101000000001010101000000000010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X30Y38, nonlinear_LMDPL
constant Tile_X30Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X31Y38, linear_LMDPL
constant Tile_X31Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000110011001100110";
--X32Y38, linear_LMDPL
constant Tile_X32Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X33Y38, nonlinear_LMDPL
constant Tile_X33Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000110011001100110011001100110011000000000000000000";
--X34Y38, linear_LMDPL
constant Tile_X34Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X35Y38, linear_LMDPL
constant Tile_X35Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X36Y38, nonlinear_LMDPL
constant Tile_X36Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000111011101110111001000100010001000000000000000000";
--X37Y38, linear_LMDPL
constant Tile_X37Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X38Y38, linear_LMDPL
constant Tile_X38Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000101010101000000000101010101010101000000000000000000000000000000000101010101010101";
--X39Y38, nonlinear_LMDPL
constant Tile_X39Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y38, linear_LMDPL
constant Tile_X40Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000101010100000000000000000101010100000000000000000000000001111111101010101101010100000000010101010000000000000000000000000000000000000000010101010000000000101010111111111000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000011001100110011";
--X41Y38, linear_LMDPL
constant Tile_X41Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000001100110011001101000100010001000000000000000000";
--X42Y38, nonlinear_LMDPL
constant Tile_X42Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101011010101000000000010101010000000010101010000000000000000000000000101010101010101000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000011001100110011";
--X43Y38, linear_LMDPL
constant Tile_X43Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000001010101000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X44Y38, linear_LMDPL
constant Tile_X44Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X45Y38, nonlinear_LMDPL
constant Tile_X45Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000000001000100010001";
--X46Y38, linear_LMDPL
constant Tile_X46Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010101010101000000000000000000101010110101010000000000000000010101010111111111010101000000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X47Y38, linear_LMDPL
constant Tile_X47Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000001010101010101010000000000000000000000000000000001010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X48Y38, nonlinear_LMDPL
constant Tile_X48Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101011111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000001010101000000000101010100000000000000000000000010101010000000000000000010101010010001000100010000000000000000000000000000000000111011101110111000100010001000100000000000000000";
--X49Y38, linear_LMDPL
constant Tile_X49Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101000000000101010100000000010101010000000000000000001010101000000001010101000000000010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X50Y38, linear_LMDPL
constant Tile_X50Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000000000000000000010101010101010101010101000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X51Y38, nonlinear_LMDPL
constant Tile_X51Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000001010101010101010000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X52Y38, linear_LMDPL
constant Tile_X52Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010111111111000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100";
--X53Y38, linear_LMDPL
constant Tile_X53Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000111111110000000000000000000000000000000000000000010101010000000000000000000000001010101000000000101010100101010100000000000000000000000000000000101010101010101000000000010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X54Y38, nonlinear_LMDPL
constant Tile_X54Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001111111100000000000000000101010110101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X55Y38, linear_LMDPL
constant Tile_X55Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011011001100110011000000000000000000";
--X56Y38, linear_LMDPL
constant Tile_X56Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X57Y38, nonlinear_LMDPL
constant Tile_X57Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101101010100000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X58Y38, linear_LMDPL
constant Tile_X58Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101010101010000000000000000011111111101010101010101011111111010001000100010000000000000000000000000000000000001000100010001000110011001100110000000000000000";
--X59Y38, linear_LMDPL
constant Tile_X59Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000100010001000100";
--X60Y38, nonlinear_LMDPL
constant Tile_X60Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000111111110000000000000000010101010000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000011101110111011110001000100010000000000000000000";
--X61Y38, linear_LMDPL
constant Tile_X61Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001100110011001100";
--X62Y38, linear_LMDPL
constant Tile_X62Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000100010001000100000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X63Y38, nonlinear_LMDPL
constant Tile_X63Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000001010101010101011010101001010101000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000010001000100010";
--X64Y38, linear_LMDPL
constant Tile_X64Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101011010101010101010000000000000000011111111101010101010101000000000010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X65Y38, linear_LMDPL
constant Tile_X65Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000001010101001010101000000000000000000000000000000000000000000000000000100010001000100000000010101010100010001000100000000000000000000000000000000000101010101010101";
--X66Y38, nonlinear_LMDPL
constant Tile_X66Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y38, linear_LMDPL
constant Tile_X67Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000000000000010101010101010101010101000000000000100010001000100000000101010100010001000100010000000000000000000000000000000001010101010101010";
--X68Y38, linear_LMDPL
constant Tile_X68Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000000000000000000000110011001100110000000000000000";
--X69Y38, nonlinear_LMDPL
constant Tile_X69Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010000000001010101010101010000100010001000100000000101010100010001000100010000000000000000000000000000000000000000000000000";
--X70Y38, linear_LMDPL
constant Tile_X70Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X71Y38, linear_LMDPL
constant Tile_X71Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010000000001010101000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000011001100110011";
--X72Y38, nonlinear_LMDPL
constant Tile_X72Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000010101010000100010001000100000000000000000101010101010101000000000000000000000000000000000100010001000100";
--X73Y38, linear_LMDPL
constant Tile_X73Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001011101110111011";
--X74Y38, linear_LMDPL
constant Tile_X74Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X75Y38, nonlinear_LMDPL
constant Tile_X75Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000001010101000000000000000000000000101010101010101000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X76Y38, linear_LMDPL
constant Tile_X76Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000001111111100000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000010101010010101010101010100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X77Y38, linear_LMDPL
constant Tile_X77Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000101010100000000000000000110011001100110000110011001100110000000000000000";
--X78Y38, ctrl_to_sec
constant Tile_X78Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y38, combined_WDDL
constant Tile_X79Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000011110000101010100000000000000000000000000101010100000000101000000000000000100010000000001001100100000000";
--X80Y38, combined_WDDL
constant Tile_X80Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y38, ctrl_IO
constant Tile_X81Y38_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y39, W_IO_custom
constant Tile_X0Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y39, linear_LMDPL
constant Tile_X1Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000011111111000000001010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X2Y39, linear_LMDPL
constant Tile_X2Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000001010101001010101000000000000000000000000000000000000000000000000010101010101010100000000010101010010001000100010000000000000000001000100010001000000000000000000";
--X3Y39, nonlinear_LMDPL
constant Tile_X3Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000010101010000000000000000000000001010101001010101000000000000000000000000010101010000000010101010010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X4Y39, linear_LMDPL
constant Tile_X4Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000001010101000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X5Y39, linear_LMDPL
constant Tile_X5Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000101010100000000101010100000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X6Y39, nonlinear_LMDPL
constant Tile_X6Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010101010101011111111010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X7Y39, linear_LMDPL
constant Tile_X7Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X8Y39, linear_LMDPL
constant Tile_X8Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X9Y39, nonlinear_LMDPL
constant Tile_X9Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X10Y39, linear_LMDPL
constant Tile_X10Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000011111111000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001110111011101110000000000000000";
--X11Y39, linear_LMDPL
constant Tile_X11Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X12Y39, nonlinear_LMDPL
constant Tile_X12Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000100010001000100000000000000001001100110011001000000000000000000000000000000001010101010101010";
--X13Y39, linear_LMDPL
constant Tile_X13Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X14Y39, linear_LMDPL
constant Tile_X14Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X15Y39, nonlinear_LMDPL
constant Tile_X15Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000101010100000000000000000101010101010101000110011001100110000000000000000";
--X16Y39, linear_LMDPL
constant Tile_X16Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000000010001000100010000000000000000000000000000000000101110111011101101010101010101010000000000000000";
--X17Y39, linear_LMDPL
constant Tile_X17Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101101010100000000000000000000000001010101010101010000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X18Y39, nonlinear_LMDPL
constant Tile_X18Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000100010001000100000000000000000000000000000000";
--X19Y39, linear_LMDPL
constant Tile_X19Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X20Y39, linear_LMDPL
constant Tile_X20Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X21Y39, nonlinear_LMDPL
constant Tile_X21Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111101010101101010101010101000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001110111011101110";
--X22Y39, linear_LMDPL
constant Tile_X22Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001110111011101110000000000000000";
--X23Y39, linear_LMDPL
constant Tile_X23Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X24Y39, nonlinear_LMDPL
constant Tile_X24Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000011001100110011001000100010001000000000000000000";
--X25Y39, linear_LMDPL
constant Tile_X25Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X26Y39, linear_LMDPL
constant Tile_X26Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101010101010000000000000000010101010111111110000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X27Y39, nonlinear_LMDPL
constant Tile_X27Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000000100010001000100";
--X28Y39, linear_LMDPL
constant Tile_X28Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111110101010101010100101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001101110111011101";
--X29Y39, linear_LMDPL
constant Tile_X29Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000010101010000000001010101000000000000000000000000010101010000000000000000000000000001000100010001000000000000000000101010101010101";
--X30Y39, nonlinear_LMDPL
constant Tile_X30Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000101010101010101";
--X31Y39, linear_LMDPL
constant Tile_X31Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000101010100000000010101010000000000000000010101010111111110000000000000000010101010101010110101010000000000000000000000000000000000000000011111111111111110000000000000000";
--X32Y39, linear_LMDPL
constant Tile_X32Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X33Y39, nonlinear_LMDPL
constant Tile_X33Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y39, linear_LMDPL
constant Tile_X34Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000011001100110011";
--X35Y39, linear_LMDPL
constant Tile_X35Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X36Y39, nonlinear_LMDPL
constant Tile_X36Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000000000000000000";
--X37Y39, linear_LMDPL
constant Tile_X37Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000111111110000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000111011101110111";
--X38Y39, linear_LMDPL
constant Tile_X38Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X39Y39, nonlinear_LMDPL
constant Tile_X39Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000111011101110111001000100010001000000000000000000";
--X40Y39, linear_LMDPL
constant Tile_X40Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010000000000101010110101010000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X41Y39, linear_LMDPL
constant Tile_X41Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X42Y39, nonlinear_LMDPL
constant Tile_X42Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111101010101010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001001100110011001";
--X43Y39, linear_LMDPL
constant Tile_X43Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111101010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000010101010101010111111111111111110000000000000000";
--X44Y39, linear_LMDPL
constant Tile_X44Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010101010101000000000101010100000000000000000000000000101010111111111010001000100010000000000000000000000000000000000110011001100110011011101110111010000000000000000";
--X45Y39, nonlinear_LMDPL
constant Tile_X45Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X46Y39, linear_LMDPL
constant Tile_X46Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010101010101000000000101010100101010111111111000000000000000000000000101010100000000000000000010001000100010010101010000000000000000000000000010001000100010010001000100010000000000000000000";
--X47Y39, linear_LMDPL
constant Tile_X47Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000001010101000000000000000001010101010101010000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000101010101010101000000000000000001000100010001000";
--X48Y39, nonlinear_LMDPL
constant Tile_X48Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010101010110101010101010100101010100000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000101010101010101000000001111111100000000000000000101010100000000010001000100010000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X49Y39, linear_LMDPL
constant Tile_X49Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000101010110101010000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X50Y39, linear_LMDPL
constant Tile_X50Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000101010101010101101010100000000000000000000000001010101000000000000000000101010100000000000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X51Y39, nonlinear_LMDPL
constant Tile_X51Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010111111111000000000000000000000000101010100000000000000000010101010000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010001000100010000000000000000001001100110011001";
--X52Y39, linear_LMDPL
constant Tile_X52Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000000000000011111111101010101010101000000000010101010101010111111111000000001010101010101010000000000000000000000000000000000000000000000000";
--X53Y39, linear_LMDPL
constant Tile_X53Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000010101011010101000000000000000000000000010101010000000001010101000000000010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X54Y39, nonlinear_LMDPL
constant Tile_X54Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010101010101000000000000000000000000000000000101010100000000000000000011101110111011100000000000000001100110011001100";
--X55Y39, linear_LMDPL
constant Tile_X55Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010101010100101010100000000101010100000000000000000000000000000000011111111010001000100010001010101010101010000000000000000000000000000000000000000000000000000000000000000";
--X56Y39, linear_LMDPL
constant Tile_X56Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000000000001010101000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X57Y39, nonlinear_LMDPL
constant Tile_X57Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000010101010000000000000000000000000111111111010101010101010000000000000000010101010101010100101010101010101010101010101010100000000010101010110011001100110000000000000000010101010101010100000000000000000";
--X58Y39, linear_LMDPL
constant Tile_X58Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100101010100000000000000001111111100000000000000000000000010101010000000001010101010101010101010100000000000000000111111110101010100000000010101010101010110101010101010100111011101110111000000000000000010101010101010100000000000000000";
--X59Y39, linear_LMDPL
constant Tile_X59Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000010101010000000000000000111111110000000000000000101010100101010111111111000000000000000010101010101010100000000010101010000100010001000110101010101010100010001000100010000000000000000000000000000000001010101010101010";
--X60Y39, nonlinear_LMDPL
constant Tile_X60Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000010101010000000000000000011001100110011011001100110011000000000000000000";
--X61Y39, linear_LMDPL
constant Tile_X61Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000011111111000100010001000100000000101010101010101010101010000000000000000000000000000000001010101010101010";
--X62Y39, linear_LMDPL
constant Tile_X62Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101001010101000000000101010110101010000000000101010111111111000100010001000100000000000000001011101110111011000000000000000000000000000000000011001100110011";
--X63Y39, nonlinear_LMDPL
constant Tile_X63Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000101010100011001100110011000000000000000000000000000000001000100010001000";
--X64Y39, linear_LMDPL
constant Tile_X64Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000100000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X65Y39, linear_LMDPL
constant Tile_X65Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111010101010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010";
--X66Y39, nonlinear_LMDPL
constant Tile_X66Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101000000000010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X67Y39, linear_LMDPL
constant Tile_X67Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001111111100000000101010100000000000000000000000001111111101010101000000000000000000000000101010100000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010101010101001010101010001000100010000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X68Y39, linear_LMDPL
constant Tile_X68Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101101010100000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X69Y39, nonlinear_LMDPL
constant Tile_X69Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000110011001100110000110011001100110000000000000000";
--X70Y39, linear_LMDPL
constant Tile_X70Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000011111111010101010000000011111111010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X71Y39, linear_LMDPL
constant Tile_X71Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X72Y39, nonlinear_LMDPL
constant Tile_X72Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101010101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X73Y39, linear_LMDPL
constant Tile_X73Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X74Y39, linear_LMDPL
constant Tile_X74Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X75Y39, nonlinear_LMDPL
constant Tile_X75Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000101010100000000001010101000000000000000010101010101010100000000010101010000100010001000100000000010101010000000000000000000000000000000000000000000000000101010101010101";
--X76Y39, linear_LMDPL
constant Tile_X76Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101011111111000000000000000000000000101010100000000010101010010101010101010100000000101010100011001100110011000000000000000010001000100010000000000000000000";
--X77Y39, linear_LMDPL
constant Tile_X77Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000100010001000100001010101010101010000000000000000";
--X78Y39, ctrl_to_sec
constant Tile_X78Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y39, combined_WDDL
constant Tile_X79Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y39, combined_WDDL
constant Tile_X80Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y39, ctrl_IO
constant Tile_X81Y39_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y40, W_IO_custom
constant Tile_X0Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y40, linear_LMDPL
constant Tile_X1Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000010101010000000000000000000000001010101011111111010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X2Y40, linear_LMDPL
constant Tile_X2Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000001010101010101010000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000100110011001100100000000000000000001000100010001";
--X3Y40, nonlinear_LMDPL
constant Tile_X3Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X4Y40, linear_LMDPL
constant Tile_X4Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100110011001100101010101010101010000000000000000";
--X5Y40, linear_LMDPL
constant Tile_X5Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X6Y40, nonlinear_LMDPL
constant Tile_X6Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X7Y40, linear_LMDPL
constant Tile_X7Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000001010101010101010000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X8Y40, linear_LMDPL
constant Tile_X8Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100000110011001100110000000000000000";
--X9Y40, nonlinear_LMDPL
constant Tile_X9Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010010001000100010000000000000000000000000000000000101110111011101110111011101110110000000000000000";
--X10Y40, linear_LMDPL
constant Tile_X10Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101010100000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X11Y40, linear_LMDPL
constant Tile_X11Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X12Y40, nonlinear_LMDPL
constant Tile_X12Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000100110011001100110101010101010100000000000000000";
--X13Y40, linear_LMDPL
constant Tile_X13Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000111111110000000000000000101010100000000000000000111111110000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X14Y40, linear_LMDPL
constant Tile_X14Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X15Y40, nonlinear_LMDPL
constant Tile_X15Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101000010001000100010000000000000000";
--X16Y40, linear_LMDPL
constant Tile_X16Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010";
--X17Y40, linear_LMDPL
constant Tile_X17Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000010101011010101000000000000000000000000011111111000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X18Y40, nonlinear_LMDPL
constant Tile_X18Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000011001100110011";
--X19Y40, linear_LMDPL
constant Tile_X19Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101110111011101100000000000000001010101010101010";
--X20Y40, linear_LMDPL
constant Tile_X20Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X21Y40, nonlinear_LMDPL
constant Tile_X21Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000101010100000000101010101010101000000000000000001010101000000000000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X22Y40, linear_LMDPL
constant Tile_X22Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000110011001100110000000000000000001011101110111011";
--X23Y40, linear_LMDPL
constant Tile_X23Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X24Y40, nonlinear_LMDPL
constant Tile_X24Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000001100110011001100000000000000001001100110011001";
--X25Y40, linear_LMDPL
constant Tile_X25Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000101010101000100010001000000000000000000011011101110111010000000000000000";
--X26Y40, linear_LMDPL
constant Tile_X26Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000010101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X27Y40, nonlinear_LMDPL
constant Tile_X27Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X28Y40, linear_LMDPL
constant Tile_X28Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000111111110000000010101010101010101010101010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X29Y40, linear_LMDPL
constant Tile_X29Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000010101010000000001010101000000000010101010101010111111111000000001010101010101010000000000000000000000000000000000000000000000000";
--X30Y40, nonlinear_LMDPL
constant Tile_X30Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000101010101010101";
--X31Y40, linear_LMDPL
constant Tile_X31Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000110011001100110";
--X32Y40, linear_LMDPL
constant Tile_X32Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X33Y40, nonlinear_LMDPL
constant Tile_X33Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y40, linear_LMDPL
constant Tile_X34Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X35Y40, linear_LMDPL
constant Tile_X35Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000000111011101110111";
--X36Y40, nonlinear_LMDPL
constant Tile_X36Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101001010101000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y40, linear_LMDPL
constant Tile_X37Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101111111111010101001010101000000000000000010101010101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X38Y40, linear_LMDPL
constant Tile_X38Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101011111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000101010101010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X39Y40, nonlinear_LMDPL
constant Tile_X39Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X40Y40, linear_LMDPL
constant Tile_X40Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000001010101010101010000000000101010110101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010001010101010101010000000000000000";
--X41Y40, linear_LMDPL
constant Tile_X41Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111111111110000000000000000010101010101010100000000101010101000100010001000000000000000000001000100010001000000000000000000";
--X42Y40, nonlinear_LMDPL
constant Tile_X42Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101011111111010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X43Y40, linear_LMDPL
constant Tile_X43Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000101010101010101010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X44Y40, linear_LMDPL
constant Tile_X44Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100101010100000000101010100101010100000000000000000000000000000000000000000101010100000000010001000100010000000000101010100000000000000000000000000000000010101010101010100000000000000000";
--X45Y40, nonlinear_LMDPL
constant Tile_X45Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101001100110011001000000000000000010001000100010000000000000000000";
--X46Y40, linear_LMDPL
constant Tile_X46Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000010101010000000001010101000000000000000000000000101010100000000000000000101010100000000010101010000000000000000010101010101010100101010111111111000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X47Y40, linear_LMDPL
constant Tile_X47Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101000000000111111111010101010101010000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X48Y40, nonlinear_LMDPL
constant Tile_X48Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000101010101010101010101010000000000000000000000001010101000000000000000001010101000000000000000001010101000000000000000001010101000000000010101010101010111111111000000001101110111011101000000000000000010011001100110010000000000000000";
--X49Y40, linear_LMDPL
constant Tile_X49Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000000000000010101010111111111010101001010101000000000000000000000000000000000000000000000000110011001100110000000000000000000100010001000100";
--X50Y40, linear_LMDPL
constant Tile_X50Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101101010101010101000000000000100010001000100000000111111110000000000000000000000000000000000000000000000001000100010001000";
--X51Y40, nonlinear_LMDPL
constant Tile_X51Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000111011101110111000000000000000000000000000000000";
--X52Y40, linear_LMDPL
constant Tile_X52Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101000000000000000001010101001010101000000000000000000000000101010100101010100000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X53Y40, linear_LMDPL
constant Tile_X53Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111010101010101010100000000000000000000000000000000101010100000000000000000010101010000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000011111111111111110000000000000000";
--X54Y40, nonlinear_LMDPL
constant Tile_X54Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000001111111100000000000000000101010110101010101010100000000000000000010101011010101000000000010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X55Y40, linear_LMDPL
constant Tile_X55Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010101010101010101000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X56Y40, linear_LMDPL
constant Tile_X56Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X57Y40, nonlinear_LMDPL
constant Tile_X57Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010101010101111111100000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000010101010000000000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X58Y40, linear_LMDPL
constant Tile_X58Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010111111111010101001010101101010100000000000000000101010100000000001010101010001000100010000000000000000000000000000000000100010001000100011011101110111010000000000000000";
--X59Y40, linear_LMDPL
constant Tile_X59Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000111111110101010100000000000000000000000000000000000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X60Y40, nonlinear_LMDPL
constant Tile_X60Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000101010101010101000000000000000000000000010101010101010100000000000100010001000100000000010101011011101110111011000000000000000000000000000000001010101010101010";
--X61Y40, linear_LMDPL
constant Tile_X61Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000001010101000000000000000001111111110101010000000000000000000000000101010100000000000000000000000001010101000000000000000001010101001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X62Y40, linear_LMDPL
constant Tile_X62Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111000000001010101010101010000000001010101000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101000000000000000000000000011111111101010101010101000000000000100010001000100000000010101010100010001000100000000000000000000000000000000001011101110111011";
--X63Y40, nonlinear_LMDPL
constant Tile_X63Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000010101010000000000000000000000001010101001010101000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000010001000100010";
--X64Y40, linear_LMDPL
constant Tile_X64Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000010101010101010100000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000101010101010101";
--X65Y40, linear_LMDPL
constant Tile_X65Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000101010100000000000100010001000100000000101010100101010101010101000000000000000000000000000000001000100010001000";
--X66Y40, nonlinear_LMDPL
constant Tile_X66Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000010101010101010100101010100000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X67Y40, linear_LMDPL
constant Tile_X67Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000011111111101010100000000000000000010001000100010000000000101010100000000000000000001000100010001011011101110111010000000000000000";
--X68Y40, linear_LMDPL
constant Tile_X68Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010010101010101010110101010000000000100010001000100000000000000000000000000000000000000000000000000";
--X69Y40, nonlinear_LMDPL
constant Tile_X69Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010000000001111111110101010010101010101010100000000101010100010001000100010000000000000000010111011101110110000000000000000";
--X70Y40, linear_LMDPL
constant Tile_X70Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X71Y40, linear_LMDPL
constant Tile_X71Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000100010001000100";
--X72Y40, nonlinear_LMDPL
constant Tile_X72Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101001010101010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X73Y40, linear_LMDPL
constant Tile_X73Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000011111111010101011010101010101010010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X74Y40, linear_LMDPL
constant Tile_X74Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111101010101000000000000000000000000101010101010101010101010010101010101010100000000000000000011001100110011000000000000000011011101110111010000000000000000";
--X75Y40, nonlinear_LMDPL
constant Tile_X75Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000000001000100010001000000000000000000000000000000000010001000100010";
--X76Y40, linear_LMDPL
constant Tile_X76Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000001001100110011001000000000000000010111011101110110000000000000000";
--X77Y40, linear_LMDPL
constant Tile_X77Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010101111111111111111000000000000000000000000000000000000000000000000";
--X78Y40, ctrl_to_sec
constant Tile_X78Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y40, combined_WDDL
constant Tile_X79Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y40, combined_WDDL
constant Tile_X80Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y40, ctrl_IO
constant Tile_X81Y40_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y41, W_IO_custom
constant Tile_X0Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y41, linear_LMDPL
constant Tile_X1Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000001010101000000000111111110000000000000000000000001010101010101010010101010101010100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X2Y41, linear_LMDPL
constant Tile_X2Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000001010101000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X3Y41, nonlinear_LMDPL
constant Tile_X3Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000100110011001100111001100110011000000000000000000";
--X4Y41, linear_LMDPL
constant Tile_X4Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X5Y41, linear_LMDPL
constant Tile_X5Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101010101010000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X6Y41, nonlinear_LMDPL
constant Tile_X6Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X7Y41, linear_LMDPL
constant Tile_X7Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000111111110000000010101010010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X8Y41, linear_LMDPL
constant Tile_X8Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X9Y41, nonlinear_LMDPL
constant Tile_X9Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X10Y41, linear_LMDPL
constant Tile_X10Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X11Y41, linear_LMDPL
constant Tile_X11Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000010101011101110111011101000000000000000000000000000000001101110111011101";
--X12Y41, nonlinear_LMDPL
constant Tile_X12Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000010101010000000000000000001000100010001000010001000100010000000000000000";
--X13Y41, linear_LMDPL
constant Tile_X13Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000001111111100000000010101010101010100000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010101010101010100000000000000000000000000000000";
--X14Y41, linear_LMDPL
constant Tile_X14Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X15Y41, nonlinear_LMDPL
constant Tile_X15Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010100110011001100110000000000000000000000000000000000011001100110011";
--X16Y41, linear_LMDPL
constant Tile_X16Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X17Y41, linear_LMDPL
constant Tile_X17Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001101110111011101";
--X18Y41, nonlinear_LMDPL
constant Tile_X18Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010101010000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X19Y41, linear_LMDPL
constant Tile_X19Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X20Y41, linear_LMDPL
constant Tile_X20Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010101010101000000000000000000011001100110011";
--X21Y41, nonlinear_LMDPL
constant Tile_X21Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100101010100000000000000001111111100000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000110011001100110";
--X22Y41, linear_LMDPL
constant Tile_X22Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X23Y41, linear_LMDPL
constant Tile_X23Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001011101110111011";
--X24Y41, nonlinear_LMDPL
constant Tile_X24Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000010001000100010000000000000000001001100110011001";
--X25Y41, linear_LMDPL
constant Tile_X25Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010101010101010111111111000000001010101010101010000000000000000011011101110111010000000000000000";
--X26Y41, linear_LMDPL
constant Tile_X26Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000010101010000000000000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X27Y41, nonlinear_LMDPL
constant Tile_X27Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X28Y41, linear_LMDPL
constant Tile_X28Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010101010101010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X29Y41, linear_LMDPL
constant Tile_X29Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010111111110000000001010101101010100000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000001010101000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X30Y41, nonlinear_LMDPL
constant Tile_X30Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X31Y41, linear_LMDPL
constant Tile_X31Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000101010101010101";
--X32Y41, linear_LMDPL
constant Tile_X32Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111011100000000000000000100010001000100";
--X33Y41, nonlinear_LMDPL
constant Tile_X33Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X34Y41, linear_LMDPL
constant Tile_X34Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010110101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X35Y41, linear_LMDPL
constant Tile_X35Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X36Y41, nonlinear_LMDPL
constant Tile_X36Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y41, linear_LMDPL
constant Tile_X37Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000101010110101010000000000000000000000000101010100000000000000000000100010001000100000000010101010100010001000100000000000000000000000000000000000111011101110111";
--X38Y41, linear_LMDPL
constant Tile_X38Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010000000000000000111111110000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000100010001000100";
--X39Y41, nonlinear_LMDPL
constant Tile_X39Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X40Y41, linear_LMDPL
constant Tile_X40Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101010101010000000000000000010101010000000000000000000000000000000000101010110101010010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X41Y41, linear_LMDPL
constant Tile_X41Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100101010111111111000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X42Y41, nonlinear_LMDPL
constant Tile_X42Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X43Y41, linear_LMDPL
constant Tile_X43Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101101010100000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000000101010101010101000000000000000000100010001000100000000000000000";
--X44Y41, linear_LMDPL
constant Tile_X44Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000101010101010101101010101010101000000000101010100000000000000000000000000000000000000000101010101010101001010101101010100000000000000000000000000101010100000000000100010001000100000000000000000101010101010101000000000000000000000000000000000010001000100010";
--X45Y41, nonlinear_LMDPL
constant Tile_X45Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001001100110011001";
--X46Y41, linear_LMDPL
constant Tile_X46Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101010101010000000000000000000000000000000000000000101010100101010101010101101010100000000010101010000000000000000001010101101010101010101001010101010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X47Y41, linear_LMDPL
constant Tile_X47Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111100000000000000001111111101010101101010100000000000000000101010100000000001010101000000000101010111111111000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X48Y41, nonlinear_LMDPL
constant Tile_X48Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000001010101000000000000000001010101000000000000000000000000000000001010101000000000101010100101010100000000000000000000000000000000000000000101010100000000010101010101010100000000000000001011101110111011000000000000000001000100010001000000000000000000";
--X49Y41, linear_LMDPL
constant Tile_X49Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000101010100000000101010101010101000000000000000000000000010101010101010101010101010101010010001000100010000000000010101010000000000000000010001000100010010001000100010000000000000000000";
--X50Y41, linear_LMDPL
constant Tile_X50Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000000000000000000000000000000101010100000000000000000000000000000000010101010000000010101010010101010000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000100010001000100011001100110011000000000000000000";
--X51Y41, nonlinear_LMDPL
constant Tile_X51Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000011111111010001000100010000000000101010100000000000000000100110011001100110111011101110110000000000000000";
--X52Y41, linear_LMDPL
constant Tile_X52Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000111111110000000000000000000000001010101000000000000000000000000010101010000000000000000000000000010101010000000000000000000000001010101000000000000000001010101000000000000000000000000010101010010101011010101000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000101010101010101";
--X53Y41, linear_LMDPL
constant Tile_X53Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010011011101110111010000000000000000";
--X54Y41, nonlinear_LMDPL
constant Tile_X54Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010101010101000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000101010100000000010101010101010100000000101010101011101110111011000000000000000011011101110111010000000000000000";
--X55Y41, linear_LMDPL
constant Tile_X55Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000101010100000000000000000010101010000000000000000000000001010101010101010101010101010101011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001001100110011001";
--X56Y41, linear_LMDPL
constant Tile_X56Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010101010000000000000000000000001010101000000000000000000000000010101010101010101010101000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X57Y41, nonlinear_LMDPL
constant Tile_X57Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000101010110101010000000000000000010101010010101010000000000000000000100010001000100000000010101011110111011101110000000000000000000000000000000000100010001000100";
--X58Y41, linear_LMDPL
constant Tile_X58Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000101010110101010000000001010101000000000101010100000000000000000000000000000000010101010000000001010101010101010000000000000000000000000111111110000000000000000010001000100010011111111101010100000000000000000010001000100010000110011001100110000000000000000";
--X59Y41, linear_LMDPL
constant Tile_X59Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000000000010101010010101010000000010101010000100010001000100000000101010100111011101110111000000000000000000000000000000000000000000000000";
--X60Y41, nonlinear_LMDPL
constant Tile_X60Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000010101011010101011111111010001000100010000000000101010100000000000000000000100010001000110001000100010000000000000000000";
--X61Y41, linear_LMDPL
constant Tile_X61Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000101010100000000010101011010101010101010000000000000000000000000010101010000000010101010000000000000000000000000101010100000000000000000100010001000100000000000000000000111011101110111";
--X62Y41, linear_LMDPL
constant Tile_X62Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010101111111100000000000000000000000001010101000000001010101000000000000000000000000000000000101010101010101010101010010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X63Y41, nonlinear_LMDPL
constant Tile_X63Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101011111111000100010001000100000000101010101100110011001100000000000000000000000000000000001001100110011001";
--X64Y41, linear_LMDPL
constant Tile_X64Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000101010100100010001000100000000000000000000000000000000000101010101010101";
--X65Y41, linear_LMDPL
constant Tile_X65Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101111111110000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000001010101011111111000100010001000100000000010101010100010001000100000000000000000000000000000000001100110011001100";
--X66Y41, nonlinear_LMDPL
constant Tile_X66Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000101010101010101";
--X67Y41, linear_LMDPL
constant Tile_X67Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000010001000100010000110011001100110000000000000000";
--X68Y41, linear_LMDPL
constant Tile_X68Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000010101010010101010101010100000000010101010101010101010101000000000000000011011101110111010000000000000000";
--X69Y41, nonlinear_LMDPL
constant Tile_X69Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X70Y41, linear_LMDPL
constant Tile_X70Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000010101010101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X71Y41, linear_LMDPL
constant Tile_X71Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X72Y41, nonlinear_LMDPL
constant Tile_X72Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000100010001000100";
--X73Y41, linear_LMDPL
constant Tile_X73Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X74Y41, linear_LMDPL
constant Tile_X74Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000010101010101010100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X75Y41, nonlinear_LMDPL
constant Tile_X75Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010101010101111111100000000010101010101010100000000010101010011001100110011000000000000000001010101010101010000000000000000";
--X76Y41, linear_LMDPL
constant Tile_X76Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000010101010000000001111111100000000000000000000000011111111000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010";
--X77Y41, linear_LMDPL
constant Tile_X77Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000001010101000000000000000000000000010101010000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000001100110011001101110111011101110000000000000000";
--X78Y41, ctrl_to_sec
constant Tile_X78Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y41, combined_WDDL
constant Tile_X79Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y41, combined_WDDL
constant Tile_X80Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y41, ctrl_IO
constant Tile_X81Y41_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y42, W_IO_custom
constant Tile_X0Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y42, linear_LMDPL
constant Tile_X1Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001011101110111011000000000000000000000000000000000001000100010001";
--X2Y42, linear_LMDPL
constant Tile_X2Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000010001000100010";
--X3Y42, nonlinear_LMDPL
constant Tile_X3Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101010101010010001000100010011111111000000000000000000000000000100010001000110001000100010000000000000000000";
--X4Y42, linear_LMDPL
constant Tile_X4Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X5Y42, linear_LMDPL
constant Tile_X5Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001010101010101010";
--X6Y42, nonlinear_LMDPL
constant Tile_X6Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X7Y42, linear_LMDPL
constant Tile_X7Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X8Y42, linear_LMDPL
constant Tile_X8Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000101110111011101100000000000000000100010001000100";
--X9Y42, nonlinear_LMDPL
constant Tile_X9Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111011101110111010000000000000000";
--X10Y42, linear_LMDPL
constant Tile_X10Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X11Y42, linear_LMDPL
constant Tile_X11Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X12Y42, nonlinear_LMDPL
constant Tile_X12Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000000000000000000";
--X13Y42, linear_LMDPL
constant Tile_X13Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X14Y42, linear_LMDPL
constant Tile_X14Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011";
--X15Y42, nonlinear_LMDPL
constant Tile_X15Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X16Y42, linear_LMDPL
constant Tile_X16Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X17Y42, linear_LMDPL
constant Tile_X17Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100";
--X18Y42, nonlinear_LMDPL
constant Tile_X18Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X19Y42, linear_LMDPL
constant Tile_X19Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000101010100000000000000000000000000000000000000000000000000010001000100010";
--X20Y42, linear_LMDPL
constant Tile_X20Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X21Y42, nonlinear_LMDPL
constant Tile_X21Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010101010101000000000111111111010101000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110010011001100110010000000000000000";
--X22Y42, linear_LMDPL
constant Tile_X22Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010111111111101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X23Y42, linear_LMDPL
constant Tile_X23Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101110111011101100000000000000000000000000000000";
--X24Y42, nonlinear_LMDPL
constant Tile_X24Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000100010001000100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X25Y42, linear_LMDPL
constant Tile_X25Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000001010101010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X26Y42, linear_LMDPL
constant Tile_X26Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X27Y42, nonlinear_LMDPL
constant Tile_X27Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X28Y42, linear_LMDPL
constant Tile_X28Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000011011101110111010000000000000000";
--X29Y42, linear_LMDPL
constant Tile_X29Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010111111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000010101010000000001010101000000000010001000100010010101010000000000000000000000000001000100010001000000000000000000000000000000000";
--X30Y42, nonlinear_LMDPL
constant Tile_X30Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000100010001000100";
--X31Y42, linear_LMDPL
constant Tile_X31Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001011111111111111110000000000000000";
--X32Y42, linear_LMDPL
constant Tile_X32Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000001100110011001111011101110111010000000000000000";
--X33Y42, nonlinear_LMDPL
constant Tile_X33Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000101010100000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X34Y42, linear_LMDPL
constant Tile_X34Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X35Y42, linear_LMDPL
constant Tile_X35Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000111011101110111";
--X36Y42, nonlinear_LMDPL
constant Tile_X36Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y42, linear_LMDPL
constant Tile_X37Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000010101010101010100000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X38Y42, linear_LMDPL
constant Tile_X38Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010101010000000000000000000000000111111110000000011111111000000000000000001010101000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X39Y42, nonlinear_LMDPL
constant Tile_X39Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000111011101110111001000100010001000000000000000000";
--X40Y42, linear_LMDPL
constant Tile_X40Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111101010100101010100000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010110101010010001000100010000000000000000000000000000000000001100110011001101110111011101110000000000000000";
--X41Y42, linear_LMDPL
constant Tile_X41Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000010101010000000000000000010101010101010100000000101010100111011101110111000000000000000011011101110111010000000000000000";
--X42Y42, nonlinear_LMDPL
constant Tile_X42Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101001010101010001000100010000000000000000000000000000000000001000100010001000010001000100010000000000000000";
--X43Y42, linear_LMDPL
constant Tile_X43Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000000000000000000001010101010101010010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X44Y42, linear_LMDPL
constant Tile_X44Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010101010101000000000101010101010101010101010101010100000000000000000000000001010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X45Y42, nonlinear_LMDPL
constant Tile_X45Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000100110011001100100100010001000100000000000000000";
--X46Y42, linear_LMDPL
constant Tile_X46Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000010101011010101000000000000000000000000000000000101010101010101011111111101010100101010110101010000000000000000010101010101010100101010100000000000100010001000110101010000000001010101010101010000000000000000000000000000000001010101010101010";
--X47Y42, linear_LMDPL
constant Tile_X47Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X48Y42, nonlinear_LMDPL
constant Tile_X48Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101010101011111111110101010000000000000000000000000000000000101010100000000010101010101010100000000000000000101010100000000000000000101010100000000000100010001000100000000000000001011101110111011000000000000000000000000000000000010001000100010";
--X49Y42, linear_LMDPL
constant Tile_X49Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000010101010000000001010101000000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X50Y42, linear_LMDPL
constant Tile_X50Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000010101010010101010000000001010101000000000000000001010101000000000101010100000000000000000000000001010101111111110101010100000000000100010001000100000000101010101000100010001000000000000000000000000000000000000100010001000100";
--X51Y42, nonlinear_LMDPL
constant Tile_X51Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000101010100000000000000001010101000000000000000000000000011111111010101010101010100000000010101010111011101110111000000000000000010101010101010100000000000000000";
--X52Y42, linear_LMDPL
constant Tile_X52Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000001010101000000000000000000101010100000000000000000000000001010101000000000000000010101010000000000000000000000000000000000101010100000000000000001010101001010101000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000011101110111011111111111111111110000000000000000";
--X53Y42, linear_LMDPL
constant Tile_X53Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000101010100000000010101010000000000000000000000001010101000000000000000001010101001010101000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X54Y42, nonlinear_LMDPL
constant Tile_X54Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000010101010101010100010001000100010000000000000000";
--X55Y42, linear_LMDPL
constant Tile_X55Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000011111111101010100000000000000000111111111010101010101010101010101010101010101010111111110000000000000000010101010000000000000000000100010001000110101010000000001000100010001000000000000000000000000000000000000100010001000100";
--X56Y42, linear_LMDPL
constant Tile_X56Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101011111111000000000000000000000000101010101010101000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000110011001100110";
--X57Y42, nonlinear_LMDPL
constant Tile_X57Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000001000100010001";
--X58Y42, linear_LMDPL
constant Tile_X58Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000010101010101010100000000101010100000000010101010000000001010101011111111101010100000000000000000000000000000000000000000010001000100010010101010010101010000000000000000000000000000000011001100110011000000000000000000";
--X59Y42, linear_LMDPL
constant Tile_X59Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000010101010010001000100010010101010000000000000000000000000101010101010101000100010001000100000000000000000";
--X60Y42, nonlinear_LMDPL
constant Tile_X60Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101011111111000000000101010100000000000000000000000000000000101010101010101000000000010001000100010000000000010101010000000000000000011101110111011110101010101010100000000000000000";
--X61Y42, linear_LMDPL
constant Tile_X61Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000100010001000111111111000000001000100010001000000000000000000000000000000000000010001000100010";
--X62Y42, linear_LMDPL
constant Tile_X62Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000010101010000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X63Y42, nonlinear_LMDPL
constant Tile_X63Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X64Y42, linear_LMDPL
constant Tile_X64Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000001010101011111111000000000000000000000000000000000000000001010101101010100000000000000000010001000100010000000000000000000000000000000000010101010101010100000000000000000000000000000000";
--X65Y42, linear_LMDPL
constant Tile_X65Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X66Y42, nonlinear_LMDPL
constant Tile_X66Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X67Y42, linear_LMDPL
constant Tile_X67Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000100010001000100";
--X68Y42, linear_LMDPL
constant Tile_X68Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000010101010101010100000000010101010010101010101010111111111000000001000100010001000000000000000000001000100010001000000000000000000";
--X69Y42, nonlinear_LMDPL
constant Tile_X69Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010001000100010000000000000000000";
--X70Y42, linear_LMDPL
constant Tile_X70Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010101010101010100000000000000000101010101010101000000000000000010101010101010100000000000000000";
--X71Y42, linear_LMDPL
constant Tile_X71Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001010101010101010000000000000000000000000000100010001000100000000101010100111011101110111000000000000000000000000000000001100110011001100";
--X72Y42, nonlinear_LMDPL
constant Tile_X72Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X73Y42, linear_LMDPL
constant Tile_X73Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000001100110011001111011101110111010000000000000000";
--X74Y42, linear_LMDPL
constant Tile_X74Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001000100010001000000000000000000000110011001100110000000000000000";
--X75Y42, nonlinear_LMDPL
constant Tile_X75Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101111111101010101010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X76Y42, linear_LMDPL
constant Tile_X76Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X77Y42, linear_LMDPL
constant Tile_X77Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X78Y42, ctrl_to_sec
constant Tile_X78Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000";
--X79Y42, combined_WDDL
constant Tile_X79Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y42, combined_WDDL
constant Tile_X80Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y42, ctrl_IO
constant Tile_X81Y42_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y43, W_IO_custom
constant Tile_X0Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y43, linear_LMDPL
constant Tile_X1Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000101010101010101";
--X2Y43, linear_LMDPL
constant Tile_X2Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X3Y43, nonlinear_LMDPL
constant Tile_X3Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000001010101010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X4Y43, linear_LMDPL
constant Tile_X4Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X5Y43, linear_LMDPL
constant Tile_X5Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X6Y43, nonlinear_LMDPL
constant Tile_X6Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X7Y43, linear_LMDPL
constant Tile_X7Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000001111111100000000000100010001000111111111000000001000100010001000000000000000000000000000000000000100010001000100";
--X8Y43, linear_LMDPL
constant Tile_X8Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X9Y43, nonlinear_LMDPL
constant Tile_X9Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y43, linear_LMDPL
constant Tile_X10Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010001010101000000000000000000000000000100010001000110111011101110110000000000000000";
--X11Y43, linear_LMDPL
constant Tile_X11Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111111111111110101010101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X12Y43, nonlinear_LMDPL
constant Tile_X12Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010100000000111111110000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000011001100110011001000100010001000000000000000000";
--X13Y43, linear_LMDPL
constant Tile_X13Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000001010101000000000000000000000000101010101111111100000000010101010000000010101010000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000010101011011101110111011000000000000000001110111011101110000000000000000";
--X14Y43, linear_LMDPL
constant Tile_X14Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001101110111011101";
--X15Y43, nonlinear_LMDPL
constant Tile_X15Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000101010100101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000010001000100010";
--X16Y43, linear_LMDPL
constant Tile_X16Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X17Y43, linear_LMDPL
constant Tile_X17Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000101010100000000000000000010101010101010100000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X18Y43, nonlinear_LMDPL
constant Tile_X18Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101011111111000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X19Y43, linear_LMDPL
constant Tile_X19Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000101010100000000101010100000000000000000000000000000000010101010010101010000000000000000000000001010101000000000000000000000000010101010010101010101010100000000000000000101010101010101000000000000000011001100110011000000000000000000";
--X20Y43, linear_LMDPL
constant Tile_X20Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000010101011010101001010101000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000011101110111011100000000000000000";
--X21Y43, nonlinear_LMDPL
constant Tile_X21Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101101010100101010100000000000000001111111100000000000000000000000010101010000000000000000000000000000000001010101001010101101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000100010001000100";
--X22Y43, linear_LMDPL
constant Tile_X22Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000010001000100010";
--X23Y43, linear_LMDPL
constant Tile_X23Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X24Y43, nonlinear_LMDPL
constant Tile_X24Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000011001100110011000000000000000000";
--X25Y43, linear_LMDPL
constant Tile_X25Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X26Y43, linear_LMDPL
constant Tile_X26Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000011001100110011";
--X27Y43, nonlinear_LMDPL
constant Tile_X27Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000111111110000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X28Y43, linear_LMDPL
constant Tile_X28Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011101110111011101010101010101010000000000000000";
--X29Y43, linear_LMDPL
constant Tile_X29Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000001010101000000000010101010101010100000000000000001101110111011101000000000000000011111111111111110000000000000000";
--X30Y43, nonlinear_LMDPL
constant Tile_X30Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000101010101010101";
--X31Y43, linear_LMDPL
constant Tile_X31Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X32Y43, linear_LMDPL
constant Tile_X32Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000001010101111111110000000000000000000000000000000000000000000000001010101010101010000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111";
--X33Y43, nonlinear_LMDPL
constant Tile_X33Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000011001100110011000000000000000000000000000000000";
--X34Y43, linear_LMDPL
constant Tile_X34Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111111111110000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X35Y43, linear_LMDPL
constant Tile_X35Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X36Y43, nonlinear_LMDPL
constant Tile_X36Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X37Y43, linear_LMDPL
constant Tile_X37Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010000000000000000010101010000000000101010100000000000000000000000001010101010001000100010000000000000000000000000000000000011001100110011011001100110011000000000000000000";
--X38Y43, linear_LMDPL
constant Tile_X38Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X39Y43, nonlinear_LMDPL
constant Tile_X39Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000100010001000100000000000000001011101110111011000000000000000000000000000000001000100010001000";
--X40Y43, linear_LMDPL
constant Tile_X40Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000100010001000100";
--X41Y43, linear_LMDPL
constant Tile_X41Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101001010101000000001010101000000000010101010000000000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X42Y43, nonlinear_LMDPL
constant Tile_X42Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X43Y43, linear_LMDPL
constant Tile_X43Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X44Y43, linear_LMDPL
constant Tile_X44Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011010101000000000101010101010101001010101000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X45Y43, nonlinear_LMDPL
constant Tile_X45Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000010001000100010000000000010101010000000000000000001000100010001010011001100110010000000000000000";
--X46Y43, linear_LMDPL
constant Tile_X46Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000010101010000000000000000101010101010101001010101101010101010101010101010000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000010101010101010101000100010001000000000000000000";
--X47Y43, linear_LMDPL
constant Tile_X47Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001010101011111111000000000101010100000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101000000000000000001010101000000000000000001010101000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000000000000000000000000000000000000";
--X48Y43, nonlinear_LMDPL
constant Tile_X48Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000010101011111111111111111000000000000000000000000000000001000100010001000";
--X49Y43, linear_LMDPL
constant Tile_X49Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000001010101000000000000000001010101000000000000000000000000000000000000000001010101000000000010101010101010100000000010101010010001000100010000000000000000011011101110111010000000000000000";
--X50Y43, linear_LMDPL
constant Tile_X50Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111101010101010101000000000010101010101010100000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X51Y43, nonlinear_LMDPL
constant Tile_X51Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000001010101001010101101010100000000000000000000000001010101000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111011101110111000000000000000000101010101010101";
--X52Y43, linear_LMDPL
constant Tile_X52Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000101010100000000000000000101010111111111000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X53Y43, linear_LMDPL
constant Tile_X53Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000000000000001010101101010100000000010101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X54Y43, nonlinear_LMDPL
constant Tile_X54Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101111111110000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010";
--X55Y43, linear_LMDPL
constant Tile_X55Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000000101010110101010010101011010101010101010000000000000000001010101111111110000000000000000010001000100010000000000101010100000000000000000110011001100110011001100110011000000000000000000";
--X56Y43, linear_LMDPL
constant Tile_X56Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010100000000000000000000000000000001010101011111111101010100101010100000000000000000000000000000000000000000101010100000000101010100000000000000000111111110000000000000000000000000101010100000000000000000000000010101010101010100000000001010101000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X57Y43, nonlinear_LMDPL
constant Tile_X57Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001010101001010101000000000000000001010101101010100000000000000000000000000000000000000000010101010000000000000000001100110011001100000000000000000000000000000000";
--X58Y43, linear_LMDPL
constant Tile_X58Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000001111111100000000000000000000000010101010101010100000000010101010010101010000000010101010111111110000000000000000111111110000000000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X59Y43, linear_LMDPL
constant Tile_X59Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010000000000000000000000000101010100000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X60Y43, nonlinear_LMDPL
constant Tile_X60Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000101010101010101000000000000100010001000100000000101010101011101110111011000000000000000000000000000000000000000000000000";
--X61Y43, linear_LMDPL
constant Tile_X61Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010001000100010000000000010101010000000000000000001100110011001100000000000000000000000000000000";
--X62Y43, linear_LMDPL
constant Tile_X62Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000001000100010001001110111011101110000000000000000";
--X63Y43, nonlinear_LMDPL
constant Tile_X63Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010101011101110111011000000000000000010001000100010000000000000000000";
--X64Y43, linear_LMDPL
constant Tile_X64Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000010001000100010001000100010001000000000000000000";
--X65Y43, linear_LMDPL
constant Tile_X65Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000001010101000000000000000010101010000000000000000010101010000000000000000010101010010001000100010000000000010101010000000000000000001000100010001001000100010001000000000000000000";
--X66Y43, nonlinear_LMDPL
constant Tile_X66Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X67Y43, linear_LMDPL
constant Tile_X67Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000010101010101010100000000000000000000000000000000000000000101010101010101011111111000000000000000000000000010101010000000000000000001100110011001100000000000000001011101110111011";
--X68Y43, linear_LMDPL
constant Tile_X68Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000101010100000000010101010000100010001000110101010101010100101010101010101000000000000000000000000000000001010101010101010";
--X69Y43, nonlinear_LMDPL
constant Tile_X69Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y43, linear_LMDPL
constant Tile_X70Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000001101110111011101000000000000000000110011001100110000000000000000";
--X71Y43, linear_LMDPL
constant Tile_X71Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000001010101010101010000000000000000";
--X72Y43, nonlinear_LMDPL
constant Tile_X72Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000010101010101010100000000010101010010001000100010000000000000000010111011101110110000000000000000";
--X73Y43, linear_LMDPL
constant Tile_X73Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111111010101000000000010101010101010100000000000000001010101010101010000000000000000000110011001100110000000000000000";
--X74Y43, linear_LMDPL
constant Tile_X74Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X75Y43, nonlinear_LMDPL
constant Tile_X75Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X76Y43, linear_LMDPL
constant Tile_X76Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X77Y43, linear_LMDPL
constant Tile_X77Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X78Y43, ctrl_to_sec
constant Tile_X78Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y43, combined_WDDL
constant Tile_X79Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000111110001000000000001001100100000000";
--X80Y43, combined_WDDL
constant Tile_X80Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y43, ctrl_IO
constant Tile_X81Y43_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y44, W_IO_custom
constant Tile_X0Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y44, linear_LMDPL
constant Tile_X1Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000001000100010001";
--X2Y44, linear_LMDPL
constant Tile_X2Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X3Y44, nonlinear_LMDPL
constant Tile_X3Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001001100110011001000000000000000000000000000000000010001000100010";
--X4Y44, linear_LMDPL
constant Tile_X4Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X5Y44, linear_LMDPL
constant Tile_X5Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000110011001100110000000000000000";
--X6Y44, nonlinear_LMDPL
constant Tile_X6Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000111111110101010100000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X7Y44, linear_LMDPL
constant Tile_X7Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000000100010001000110011001100110010000000000000000";
--X8Y44, linear_LMDPL
constant Tile_X8Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000111011101110111";
--X9Y44, nonlinear_LMDPL
constant Tile_X9Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y44, linear_LMDPL
constant Tile_X10Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X11Y44, linear_LMDPL
constant Tile_X11Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X12Y44, nonlinear_LMDPL
constant Tile_X12Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010101010000000000000000001010101000000000000000000000000111111110000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000001000100010001";
--X13Y44, linear_LMDPL
constant Tile_X13Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001010101010101010000000000000000";
--X14Y44, linear_LMDPL
constant Tile_X14Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000011111111000000000000000010101010000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X15Y44, nonlinear_LMDPL
constant Tile_X15Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X16Y44, linear_LMDPL
constant Tile_X16Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000100010001000100";
--X17Y44, linear_LMDPL
constant Tile_X17Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001101110111011101000000000000000000100010001000100000000000000000";
--X18Y44, nonlinear_LMDPL
constant Tile_X18Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111000000000000000000000000000000000";
--X19Y44, linear_LMDPL
constant Tile_X19Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X20Y44, linear_LMDPL
constant Tile_X20Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X21Y44, nonlinear_LMDPL
constant Tile_X21Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000101010100000000000000000000000000000000001010101000000000000000010101010111111110000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000010101010101010100000000010101011110111011101110000000000000000001000100010001000000000000000000";
--X22Y44, linear_LMDPL
constant Tile_X22Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X23Y44, linear_LMDPL
constant Tile_X23Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X24Y44, nonlinear_LMDPL
constant Tile_X24Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111011101110111000000000000000001100110011001100";
--X25Y44, linear_LMDPL
constant Tile_X25Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000000000000000100010001000100000000000000001111111111111111000000000000000000000000000000001010101010101010";
--X26Y44, linear_LMDPL
constant Tile_X26Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X27Y44, nonlinear_LMDPL
constant Tile_X27Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X28Y44, linear_LMDPL
constant Tile_X28Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X29Y44, linear_LMDPL
constant Tile_X29Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000001010101000000000010001000100010000000000000000000000000000000000101110111011101101110111011101110000000000000000";
--X30Y44, nonlinear_LMDPL
constant Tile_X30Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000010101010000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000011001100110011";
--X31Y44, linear_LMDPL
constant Tile_X31Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001110111011101110";
--X32Y44, linear_LMDPL
constant Tile_X32Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000011111111000100010001000100000000000000000100010001000100000000000000000000000000000000000110011001100110";
--X33Y44, nonlinear_LMDPL
constant Tile_X33Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111001000100010001000000000000000000";
--X34Y44, linear_LMDPL
constant Tile_X34Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000011111111000000000000000001010101101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000001010101010101010";
--X35Y44, linear_LMDPL
constant Tile_X35Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001110111011101110";
--X36Y44, nonlinear_LMDPL
constant Tile_X36Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X37Y44, linear_LMDPL
constant Tile_X37Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000010101010000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000110011001100110";
--X38Y44, linear_LMDPL
constant Tile_X38Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010110101010000000000000000011111111000000000000000010101010010001000100010010101010000000000000000000000000010001000100010011001100110011000000000000000000";
--X39Y44, nonlinear_LMDPL
constant Tile_X39Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y44, linear_LMDPL
constant Tile_X40Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X41Y44, linear_LMDPL
constant Tile_X41Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000111111110000000010101010010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000010101010101010100000000101010100000000000000000000000000000000011001100110011000000000000000000";
--X42Y44, nonlinear_LMDPL
constant Tile_X42Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000111011101110111010101010101010100000000000000000";
--X43Y44, linear_LMDPL
constant Tile_X43Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000001010101001010101000100010001000100000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X44Y44, linear_LMDPL
constant Tile_X44Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010101111111100000000101010100101010100000000101010101010101001010101101010100000000000000000000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000000101010101010101";
--X45Y44, nonlinear_LMDPL
constant Tile_X45Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000001010101000000000000000001010101010101010000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000101110111011101101000100010001000000000000000000";
--X46Y44, linear_LMDPL
constant Tile_X46Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000101010101010101010101010000000000000000000000000000000000000000011111111000100010001000111111111000000001101110111011101000000000000000000000000000000000010001000100010";
--X47Y44, linear_LMDPL
constant Tile_X47Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000101010111111111000000000000000011111111000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001000100010001000";
--X48Y44, nonlinear_LMDPL
constant Tile_X48Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X49Y44, linear_LMDPL
constant Tile_X49Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000101010100000000101010101010101000000000000000000000000001010101101010101010101011111111000100010001000100000000111111111101110111011101000000000000000000000000000000000100010001000100";
--X50Y44, linear_LMDPL
constant Tile_X50Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010111111111000000001010101000000000000000001010101000000000010001000100010000000000101010100000000000000000100010001000100011101110111011100000000000000000";
--X51Y44, nonlinear_LMDPL
constant Tile_X51Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000010101010000000000000000000000001010101000000000000000001010101000000000000000001010101011111111010101010000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000001000100010001";
--X52Y44, linear_LMDPL
constant Tile_X52Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000010101010010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000001000100010001000000000000000000";
--X53Y44, linear_LMDPL
constant Tile_X53Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101010101010000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000001010101000000000000000010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X54Y44, nonlinear_LMDPL
constant Tile_X54Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X55Y44, linear_LMDPL
constant Tile_X55Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011111111010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010000000000101010110101010000000000000000000000000101010100000000011111111010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X56Y44, linear_LMDPL
constant Tile_X56Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X57Y44, nonlinear_LMDPL
constant Tile_X57Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000010001000100010";
--X58Y44, linear_LMDPL
constant Tile_X58Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000010101010101010100000000010101010111111111010101010101010000000000000000000000000111111110000000000000000010001000100010010101010010101010000000000000000000000000000000011001100110011000000000000000000";
--X59Y44, linear_LMDPL
constant Tile_X59Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000111111110000000010101010101010101010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100101010100000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X60Y44, nonlinear_LMDPL
constant Tile_X60Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000010101010000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111011001100110011000000000000000000";
--X61Y44, linear_LMDPL
constant Tile_X61Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010001000100010000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X62Y44, linear_LMDPL
constant Tile_X62Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000010101010000000000000000001100110011001100110011001100110000000000000000";
--X63Y44, nonlinear_LMDPL
constant Tile_X63Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X64Y44, linear_LMDPL
constant Tile_X64Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000101010100000000011111111000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X65Y44, linear_LMDPL
constant Tile_X65Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010101010101010100000000000000000000000000000000";
--X66Y44, nonlinear_LMDPL
constant Tile_X66Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y44, linear_LMDPL
constant Tile_X67Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000000111011101110111000000000000000001000100010001000000000000000000";
--X68Y44, linear_LMDPL
constant Tile_X68Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000010101010010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X69Y44, nonlinear_LMDPL
constant Tile_X69Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y44, linear_LMDPL
constant Tile_X70Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X71Y44, linear_LMDPL
constant Tile_X71Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000001010101010101010000000000000000000000000010101010101010100000000101010100100010001000100000000000000000000110011001100110000000000000000";
--X72Y44, nonlinear_LMDPL
constant Tile_X72Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X73Y44, linear_LMDPL
constant Tile_X73Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000001100110011001110111011101110110000000000000000";
--X74Y44, linear_LMDPL
constant Tile_X74Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X75Y44, nonlinear_LMDPL
constant Tile_X75Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X76Y44, linear_LMDPL
constant Tile_X76Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X77Y44, linear_LMDPL
constant Tile_X77Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110111011101110110000000000000000";
--X78Y44, ctrl_to_sec
constant Tile_X78Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y44, combined_WDDL
constant Tile_X79Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y44, combined_WDDL
constant Tile_X80Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y44, ctrl_IO
constant Tile_X81Y44_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y45, W_IO_custom
constant Tile_X0Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y45, linear_LMDPL
constant Tile_X1Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000111011101110111";
--X2Y45, linear_LMDPL
constant Tile_X2Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X3Y45, nonlinear_LMDPL
constant Tile_X3Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X4Y45, linear_LMDPL
constant Tile_X4Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000100010001000100000000010101010100010001000100000000000000000000000000000000000000000000000000";
--X5Y45, linear_LMDPL
constant Tile_X5Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X6Y45, nonlinear_LMDPL
constant Tile_X6Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000000100010001000110011001100110010000000000000000";
--X7Y45, linear_LMDPL
constant Tile_X7Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X8Y45, linear_LMDPL
constant Tile_X8Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000000100010001000111001100110011000000000000000000";
--X9Y45, nonlinear_LMDPL
constant Tile_X9Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001010101000000000000000000000000000000000000000000101010100000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000010001000100010";
--X10Y45, linear_LMDPL
constant Tile_X10Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X11Y45, linear_LMDPL
constant Tile_X11Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100101010101010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001110111011101110110000000000000000";
--X12Y45, nonlinear_LMDPL
constant Tile_X12Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X13Y45, linear_LMDPL
constant Tile_X13Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000011001100110011";
--X14Y45, linear_LMDPL
constant Tile_X14Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000001000100010001000000000000000000000000000000000000101010101010101";
--X15Y45, nonlinear_LMDPL
constant Tile_X15Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001001100110011001000000000000000011001100110011000000000000000000";
--X16Y45, linear_LMDPL
constant Tile_X16Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010110101010111111110000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000100010001000100";
--X17Y45, linear_LMDPL
constant Tile_X17Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X18Y45, nonlinear_LMDPL
constant Tile_X18Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111011101110111000000000000000000100010001000100";
--X19Y45, linear_LMDPL
constant Tile_X19Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010111111110101010100000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X20Y45, linear_LMDPL
constant Tile_X20Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010101111111100000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X21Y45, nonlinear_LMDPL
constant Tile_X21Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111110101010000000000000000000000000000000001010101000000000101010101010101000000000000000001010101000000000000000000000000000000000010101010101010100000000010101010011001100110011000000000000000000000000000000000000000000000000";
--X22Y45, linear_LMDPL
constant Tile_X22Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001110111011101110000000000000000";
--X23Y45, linear_LMDPL
constant Tile_X23Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X24Y45, nonlinear_LMDPL
constant Tile_X24Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000100010001000100001000100010001000000000000000000";
--X25Y45, linear_LMDPL
constant Tile_X25Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000000000000000000000000000000000000";
--X26Y45, linear_LMDPL
constant Tile_X26Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X27Y45, nonlinear_LMDPL
constant Tile_X27Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000001000100010001";
--X28Y45, linear_LMDPL
constant Tile_X28Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000101010101010101";
--X29Y45, linear_LMDPL
constant Tile_X29Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000100010001000110101010000000000000000000000000000000000000000000000000000000000011001100110011";
--X30Y45, nonlinear_LMDPL
constant Tile_X30Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000111011101110111";
--X31Y45, linear_LMDPL
constant Tile_X31Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001100110011001100";
--X32Y45, linear_LMDPL
constant Tile_X32Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000111111111010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110111011101110111010000000000000000";
--X33Y45, nonlinear_LMDPL
constant Tile_X33Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111010101010101010100000000000000000";
--X34Y45, linear_LMDPL
constant Tile_X34Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010000000000000000000000000010101010000000011111111000000000000000000000000000000000000000001010101101010101111111100000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X35Y45, linear_LMDPL
constant Tile_X35Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001110111011101110000000000000000";
--X36Y45, nonlinear_LMDPL
constant Tile_X36Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000100010001000100000000101010100110011001100110000000000000000000000000000000000100010001000100";
--X37Y45, linear_LMDPL
constant Tile_X37Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X38Y45, linear_LMDPL
constant Tile_X38Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101011010101010101010000000000000000000000000111111110000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000101010101010101";
--X39Y45, nonlinear_LMDPL
constant Tile_X39Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y45, linear_LMDPL
constant Tile_X40Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X41Y45, linear_LMDPL
constant Tile_X41Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000101010100000000010001000100010000000000111111110000000000000000001000100010001010101010101010100000000000000000";
--X42Y45, nonlinear_LMDPL
constant Tile_X42Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000001010101001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X43Y45, linear_LMDPL
constant Tile_X43Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000000101010101010101000000000000000011001100110011000000000000000000";
--X44Y45, linear_LMDPL
constant Tile_X44Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010100101010100000000101010101010101000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010101010101010110001000100010000000000000000000";
--X45Y45, nonlinear_LMDPL
constant Tile_X45Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010111111110000000000000000000000001010101001010101000000000101010110101010000000000000000000000000010101010000000000000000000100010001000100000000101010101101110111011101000000000000000000000000000000001000100010001000";
--X46Y45, linear_LMDPL
constant Tile_X46Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100101010110101010000000000000000000000000000000000000000010101010000100010001000100000000000000001111111111111111000000000000000000000000000000000111011101110111";
--X47Y45, linear_LMDPL
constant Tile_X47Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000010101010000000000000000000000000000000001010101010101010000000000101010100000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X48Y45, nonlinear_LMDPL
constant Tile_X48Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010101010101000000000010001000100010000000000101010100000000000000000101110111011101101000100010001000000000000000000";
--X49Y45, linear_LMDPL
constant Tile_X49Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000101010100000000000000000000000010101010000000001010101000000000010101011010101000000000000000000000000001010101101010101010101000000000010001000100010000000000010101010000000000000000001100110011001101000100010001000000000000000000";
--X50Y45, linear_LMDPL
constant Tile_X50Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000010101010111111110000000000000000101010100101010100000000000000000000000011111111000000000101010101010101010101010000000000000000000000000000000000000000000000000000000010101010000000000000000010101010010101011010101001010101010001000100010000000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X51Y45, nonlinear_LMDPL
constant Tile_X51Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000101010100000000000000001010101000000000111111110000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000001000100010001";
--X52Y45, linear_LMDPL
constant Tile_X52Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000001010101101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000000101010101010101";
--X53Y45, linear_LMDPL
constant Tile_X53Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000101010100101010100000000000000000000000000000000000000000000000010101010010101010101010100000000010101011101110111011101000000000000000010001000100010000000000000000000";
--X54Y45, nonlinear_LMDPL
constant Tile_X54Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000000000000000000";
--X55Y45, linear_LMDPL
constant Tile_X55Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010101010000000000000000000000000010101011010101001010101000000000000000000000000000000001111111100000000000000001111111110101010000000001010101010101010000000000000000001010101010101010000000000000000010001000100010010101010101010100000000000000000001000100010001011001100110011000000000000000000";
--X56Y45, linear_LMDPL
constant Tile_X56Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000001000100010001000000000000000000";
--X57Y45, nonlinear_LMDPL
constant Tile_X57Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000001010101000000000000000000000000000000000010101010000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000000000000000000";
--X58Y45, linear_LMDPL
constant Tile_X58Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000001111111100000000010101010000000000000000010101010000000010101010000000001010101010101010111111110000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111111111111111110000000000000000";
--X59Y45, linear_LMDPL
constant Tile_X59Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000101010100101010100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000011111111111111110000000000000000";
--X60Y45, nonlinear_LMDPL
constant Tile_X60Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000001010101000000000000000001010101000000000000000000000000000000000010101010000000010101010000100010001000100000000101010101110111011101110000000000000000000000000000000000011001100110011";
--X61Y45, linear_LMDPL
constant Tile_X61Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111111111110000000010101010000100010001000110101010101010100010001000100010000000000000000000000000000000000100010001000100";
--X62Y45, linear_LMDPL
constant Tile_X62Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000010101010100010001000100000000000000000000000000000000000100010001000100";
--X63Y45, nonlinear_LMDPL
constant Tile_X63Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110000000000000000000000000000000000011001100110011";
--X64Y45, linear_LMDPL
constant Tile_X64Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111100000000101010100000000010101010000000000000000000000000101010100000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X65Y45, linear_LMDPL
constant Tile_X65Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000010101010000000000000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000010001000100010";
--X66Y45, nonlinear_LMDPL
constant Tile_X66Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X67Y45, linear_LMDPL
constant Tile_X67Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000101010101010101010101010000000000000000000110011001100110000000000000000";
--X68Y45, linear_LMDPL
constant Tile_X68Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000000111011101110111000000000000000011111111111111110000000000000000";
--X69Y45, nonlinear_LMDPL
constant Tile_X69Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y45, linear_LMDPL
constant Tile_X70Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000100110011001100100100010001000100000000000000000";
--X71Y45, linear_LMDPL
constant Tile_X71Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X72Y45, nonlinear_LMDPL
constant Tile_X72Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X73Y45, linear_LMDPL
constant Tile_X73Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X74Y45, linear_LMDPL
constant Tile_X74Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000100010001000100001010101010101010000000000000000";
--X75Y45, nonlinear_LMDPL
constant Tile_X75Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X76Y45, linear_LMDPL
constant Tile_X76Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X77Y45, linear_LMDPL
constant Tile_X77Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X78Y45, ctrl_to_sec
constant Tile_X78Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y45, combined_WDDL
constant Tile_X79Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y45, combined_WDDL
constant Tile_X80Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y45, ctrl_IO
constant Tile_X81Y45_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y46, W_IO_custom
constant Tile_X0Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y46, linear_LMDPL
constant Tile_X1Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000010101010101010100000000000000000111011101110111000000000000000000100010001000100000000000000000";
--X2Y46, linear_LMDPL
constant Tile_X2Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X3Y46, nonlinear_LMDPL
constant Tile_X3Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X4Y46, linear_LMDPL
constant Tile_X4Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X5Y46, linear_LMDPL
constant Tile_X5Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X6Y46, nonlinear_LMDPL
constant Tile_X6Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110111011101110110000000000000000";
--X7Y46, linear_LMDPL
constant Tile_X7Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000110111011101110100000000000000000100010001000100";
--X8Y46, linear_LMDPL
constant Tile_X8Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000011101110111011100000000000000000011001100110011";
--X9Y46, nonlinear_LMDPL
constant Tile_X9Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000100010001000100000000000000000001000100010001000000000000000000000000000000000000000000000000";
--X10Y46, linear_LMDPL
constant Tile_X10Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111110101010010101010101010100000000000000001001100110011001000000000000000000100010001000100000000000000000";
--X11Y46, linear_LMDPL
constant Tile_X11Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000010101010111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001110111011101110";
--X12Y46, nonlinear_LMDPL
constant Tile_X12Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000001010101000000000000000001010101000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X13Y46, linear_LMDPL
constant Tile_X13Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000111011101110111000000000000000000110011001100110";
--X14Y46, linear_LMDPL
constant Tile_X14Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000010101010000000001111111100000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X15Y46, nonlinear_LMDPL
constant Tile_X15Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010101010000000000000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000101110111011101110011001100110010000000000000000";
--X16Y46, linear_LMDPL
constant Tile_X16Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X17Y46, linear_LMDPL
constant Tile_X17Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000100010001000100000000000000001010101010101010";
--X18Y46, nonlinear_LMDPL
constant Tile_X18Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010010001000100010000000000010101010000000000000000010101010101010100010001000100010000000000000000";
--X19Y46, linear_LMDPL
constant Tile_X19Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101010101010111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111111111111";
--X20Y46, linear_LMDPL
constant Tile_X20Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000000000000111111110000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X21Y46, nonlinear_LMDPL
constant Tile_X21Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000000100010001000100000000101010101001100110011001000000000000000000000000000000000000000000000000";
--X22Y46, linear_LMDPL
constant Tile_X22Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101110111011101100000000000000001010101010101010";
--X23Y46, linear_LMDPL
constant Tile_X23Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000001111111100000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X24Y46, nonlinear_LMDPL
constant Tile_X24Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000010101010000000001010101000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000111011101110111";
--X25Y46, linear_LMDPL
constant Tile_X25Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000001010101000000000000000001010101000000000000000011111111010101010101010100000000000000000101010101010101000000000000000000000000000000000000000000000000";
--X26Y46, linear_LMDPL
constant Tile_X26Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X27Y46, nonlinear_LMDPL
constant Tile_X27Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X28Y46, linear_LMDPL
constant Tile_X28Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111111111110000000000000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X29Y46, linear_LMDPL
constant Tile_X29Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111111010101000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000";
--X30Y46, nonlinear_LMDPL
constant Tile_X30Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000011001100110011000000000000000001010101010101010000000000000000";
--X31Y46, linear_LMDPL
constant Tile_X31Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X32Y46, linear_LMDPL
constant Tile_X32Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X33Y46, nonlinear_LMDPL
constant Tile_X33Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000011111111000000000000000000000000010101010000000000000000110011001100110000000000000000001101110111011101";
--X34Y46, linear_LMDPL
constant Tile_X34Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110001110111011101110000000000000000";
--X35Y46, linear_LMDPL
constant Tile_X35Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X36Y46, nonlinear_LMDPL
constant Tile_X36Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X37Y46, linear_LMDPL
constant Tile_X37Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010110101010000000000000000001010101101010100000000000000000010001000100010000000000000000000000000000000000001000100010001011111111111111110000000000000000";
--X38Y46, linear_LMDPL
constant Tile_X38Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101001010101000000000000000010101010101010100000000010101010010101010101010100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X39Y46, nonlinear_LMDPL
constant Tile_X39Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y46, linear_LMDPL
constant Tile_X40Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000000101010101010101000000000000000000000000000000000100010001000100";
--X41Y46, linear_LMDPL
constant Tile_X41Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010101100110011001100000000000000000000000000000000000000000000000000";
--X42Y46, nonlinear_LMDPL
constant Tile_X42Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000110011001100110000000000000000000000000000000000100010001000100";
--X43Y46, linear_LMDPL
constant Tile_X43Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110101010101010101010101010101010100000000111111110000000000000000000000000000000010001000100010000000000000000000";
--X44Y46, linear_LMDPL
constant Tile_X44Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000101010101010101000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000001111111111111111";
--X45Y46, nonlinear_LMDPL
constant Tile_X45Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000000100010001000111001100110011000000000000000000";
--X46Y46, linear_LMDPL
constant Tile_X46Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000101010101010101010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110001000100010001000000000000000000";
--X47Y46, linear_LMDPL
constant Tile_X47Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000101010100000000000000001010101010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X48Y46, nonlinear_LMDPL
constant Tile_X48Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010111111110000000000000000000000000000000001010101010101010101010100000000000000000000000000000000101010100101010100000000010101010101010100000000000000001011101110111011000000000000000001010101010101010000000000000000";
--X49Y46, linear_LMDPL
constant Tile_X49Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100101010100000000000000000000000000000000010101010101010100000000010101010000000011111111000000000000000011111111101010100101010110101010000000000000000000000000101010100000000000000000100010001000100000000000000000000110011001100110";
--X50Y46, linear_LMDPL
constant Tile_X50Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100101010100000000101010100000000000000000000000000000000000000000010101010000000010101010000000001010101000000000000000000000000010101010010101010101010100000000000000001100110011001100000000000000000011101110111011100000000000000000";
--X51Y46, nonlinear_LMDPL
constant Tile_X51Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000001010101000000000101010100000000000000000010101010101010100000000101010101101110111011101000000000000000001110111011101110000000000000000";
--X52Y46, linear_LMDPL
constant Tile_X52Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X53Y46, linear_LMDPL
constant Tile_X53Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101001010101000000000000000000000000010101010000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001100110011001100";
--X54Y46, nonlinear_LMDPL
constant Tile_X54Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000001010101010101010000000000000000";
--X55Y46, linear_LMDPL
constant Tile_X55Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000101010101010101000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110111011101110100000000000000001010101010101010";
--X56Y46, linear_LMDPL
constant Tile_X56Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X57Y46, nonlinear_LMDPL
constant Tile_X57Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X58Y46, linear_LMDPL
constant Tile_X58Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000101010100000000000000000010101010000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000010001000100010";
--X59Y46, linear_LMDPL
constant Tile_X59Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000111111110000000000000000000100010001000111111111000000001100110011001100000000000000000000000000000000000000000000000000";
--X60Y46, nonlinear_LMDPL
constant Tile_X60Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000000000001010101000000000101010100000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000001000100010001";
--X61Y46, linear_LMDPL
constant Tile_X61Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000100010001000100000000000000001000100010001000000000000000000000000000000000000111011101110111";
--X62Y46, linear_LMDPL
constant Tile_X62Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000001010101010101010";
--X63Y46, nonlinear_LMDPL
constant Tile_X63Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X64Y46, linear_LMDPL
constant Tile_X64Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X65Y46, linear_LMDPL
constant Tile_X65Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X66Y46, nonlinear_LMDPL
constant Tile_X66Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y46, linear_LMDPL
constant Tile_X67Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X68Y46, linear_LMDPL
constant Tile_X68Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010010001000100010010101010000000000000000000000000001000100010001000110011001100110000000000000000";
--X69Y46, nonlinear_LMDPL
constant Tile_X69Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X70Y46, linear_LMDPL
constant Tile_X70Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001000100010001000";
--X71Y46, linear_LMDPL
constant Tile_X71Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001011101110111011";
--X72Y46, nonlinear_LMDPL
constant Tile_X72Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X73Y46, linear_LMDPL
constant Tile_X73Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001001100110011001";
--X74Y46, linear_LMDPL
constant Tile_X74Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101";
--X75Y46, nonlinear_LMDPL
constant Tile_X75Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X76Y46, linear_LMDPL
constant Tile_X76Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110111011101110100000000000000001011101110111011";
--X77Y46, linear_LMDPL
constant Tile_X77Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000";
--X78Y46, ctrl_to_sec
constant Tile_X78Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y46, combined_WDDL
constant Tile_X79Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y46, combined_WDDL
constant Tile_X80Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y46, ctrl_IO
constant Tile_X81Y46_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y47, W_IO_custom
constant Tile_X0Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y47, linear_LMDPL
constant Tile_X1Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000001111111100000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X2Y47, linear_LMDPL
constant Tile_X2Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000000000000010101010101010100000000010101011000100010001000000000000000000010101010101010100000000000000000";
--X3Y47, nonlinear_LMDPL
constant Tile_X3Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X4Y47, linear_LMDPL
constant Tile_X4Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101010101010101010100000000111111111010101010101010000000000000000000100010001000100000000000000000";
--X5Y47, linear_LMDPL
constant Tile_X5Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X6Y47, nonlinear_LMDPL
constant Tile_X6Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101110111011101100000000000000000000000000000000";
--X7Y47, linear_LMDPL
constant Tile_X7Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001110111011101110";
--X8Y47, linear_LMDPL
constant Tile_X8Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X9Y47, nonlinear_LMDPL
constant Tile_X9Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000101010100000000000000000010101010000000000000000111111110000000010101010000000000000000010101010000000000000000001010101010001000100010000000000000000000000000000000000101010101010101010111011101110110000000000000000";
--X10Y47, linear_LMDPL
constant Tile_X10Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001011101110111011000000000000000000000000000000001011101110111011";
--X11Y47, linear_LMDPL
constant Tile_X11Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X12Y47, nonlinear_LMDPL
constant Tile_X12Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101111111100000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001011101110111011";
--X13Y47, linear_LMDPL
constant Tile_X13Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011111111110101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000010101010000000010101010010001000100010000000000101010100000000000000000001100110011001101110111011101110000000000000000";
--X14Y47, linear_LMDPL
constant Tile_X14Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010100000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101011111111000000000000000010101010000000000000000000000000010101010000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X15Y47, nonlinear_LMDPL
constant Tile_X15Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000000011001100110011";
--X16Y47, linear_LMDPL
constant Tile_X16Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X17Y47, linear_LMDPL
constant Tile_X17Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X18Y47, nonlinear_LMDPL
constant Tile_X18Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000101010100000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000001011101110111011";
--X19Y47, linear_LMDPL
constant Tile_X19Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010101010100101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X20Y47, linear_LMDPL
constant Tile_X20Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X21Y47, nonlinear_LMDPL
constant Tile_X21Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101111111110000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000111111111111111100000000000000001011101110111011";
--X22Y47, linear_LMDPL
constant Tile_X22Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111010101010101010100000000000000000000000001010101000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X23Y47, linear_LMDPL
constant Tile_X23Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001111111110101010010001000100010000000000000000000000000000000000101110111011101101000100010001000000000000000000";
--X24Y47, nonlinear_LMDPL
constant Tile_X24Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000001111111111111111000000000000000001010101000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110011001100110000100010001000100000000000000000";
--X25Y47, linear_LMDPL
constant Tile_X25Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000010101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X26Y47, linear_LMDPL
constant Tile_X26Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010101010101010101111111110101010101010101000000000000000010001000100010000000000000000000";
--X27Y47, nonlinear_LMDPL
constant Tile_X27Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110";
--X28Y47, linear_LMDPL
constant Tile_X28Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000101110111011101100000000000000001101110111011101";
--X29Y47, linear_LMDPL
constant Tile_X29Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000010101010101010101010101000000001011101110111011000000000000000010001000100010000000000000000000";
--X30Y47, nonlinear_LMDPL
constant Tile_X30Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X31Y47, linear_LMDPL
constant Tile_X31Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X32Y47, linear_LMDPL
constant Tile_X32Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001010101010101010";
--X33Y47, nonlinear_LMDPL
constant Tile_X33Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000001010101000000000000000001010101000000000000000001010101000000000010101010000000000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X34Y47, linear_LMDPL
constant Tile_X34Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X35Y47, linear_LMDPL
constant Tile_X35Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010001110111011101110000000000000000";
--X36Y47, nonlinear_LMDPL
constant Tile_X36Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000011111111010001000100010000000000101010100000000000000000101010101010101000100010001000100000000000000000";
--X37Y47, linear_LMDPL
constant Tile_X37Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X38Y47, linear_LMDPL
constant Tile_X38Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000001010101011111111101010100000000010101010010101010101010110101010000000001000100010001000000000000000000011011101110111010000000000000000";
--X39Y47, nonlinear_LMDPL
constant Tile_X39Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y47, linear_LMDPL
constant Tile_X40Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111101010100000000010101010010101010101010100000000101010101000100010001000000000000000000010101010101010100000000000000000";
--X41Y47, linear_LMDPL
constant Tile_X41Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X42Y47, nonlinear_LMDPL
constant Tile_X42Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X43Y47, linear_LMDPL
constant Tile_X43Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010101010101001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X44Y47, linear_LMDPL
constant Tile_X44Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000101010100000000000000000101010100000000000000000101010101010101000000000111111110000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X45Y47, nonlinear_LMDPL
constant Tile_X45Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000101010100000000000000001010101011111111000000000000000000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000000010001000100010000000000000000";
--X46Y47, linear_LMDPL
constant Tile_X46Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000010101010000000010101010000000000000000001010101000000000000000000000000000000000000000000000000101010100101010100000000101010100101010110101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X47Y47, linear_LMDPL
constant Tile_X47Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000101010101111111100000000000000000000000001010101000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001011101110111011";
--X48Y47, nonlinear_LMDPL
constant Tile_X48Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000010101010000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000111011101110111000000000000000000101010101010101";
--X49Y47, linear_LMDPL
constant Tile_X49Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000011111111101010101111111110101010000100010001000100000000000000001101110111011101000000000000000000000000000000000100010001000100";
--X50Y47, linear_LMDPL
constant Tile_X50Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000111111110000000000000000010101010101010100000000000000000100010001000100000000000000000011011101110111010000000000000000";
--X51Y47, nonlinear_LMDPL
constant Tile_X51Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000001010101001010101010101010000000011111111000100010001000100000000010101011100110011001100000000000000000000000000000000001000100010001000";
--X52Y47, linear_LMDPL
constant Tile_X52Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000101010100000000000000000101010101010101000000000000000000000000010101011111111110101010000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X53Y47, linear_LMDPL
constant Tile_X53Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111011101110111000000000000000001100110011001100";
--X54Y47, nonlinear_LMDPL
constant Tile_X54Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X55Y47, linear_LMDPL
constant Tile_X55Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001110111011101110";
--X56Y47, linear_LMDPL
constant Tile_X56Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X57Y47, nonlinear_LMDPL
constant Tile_X57Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111101010100000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011000110011001100110000000000000000";
--X58Y47, linear_LMDPL
constant Tile_X58Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111111111111111110000000000000000";
--X59Y47, linear_LMDPL
constant Tile_X59Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000001010101101010100000000011111111010101010101010100000000010101010100010001000100000000000000000011101110111011100000000000000000";
--X60Y47, nonlinear_LMDPL
constant Tile_X60Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001011101110111011";
--X61Y47, linear_LMDPL
constant Tile_X61Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000000000000000000000000010101010000000000000000110011001100110000000000000000001011101110111011";
--X62Y47, linear_LMDPL
constant Tile_X62Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111111010101000000000010101010000000000000000000000000000000000000000101010100000000010101010010001000100010000000000101010100000000000000000110011001100110000000000000000000000000000000000";
--X63Y47, nonlinear_LMDPL
constant Tile_X63Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X64Y47, linear_LMDPL
constant Tile_X64Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110111011101110100000000000000001000100010001000";
--X65Y47, linear_LMDPL
constant Tile_X65Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000010101010000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000111011101110111000000000000000000000000000000000";
--X66Y47, nonlinear_LMDPL
constant Tile_X66Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X67Y47, linear_LMDPL
constant Tile_X67Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X68Y47, linear_LMDPL
constant Tile_X68Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000100010001000111111111000000000101010101010101000000000000000000000000000000001101110111011101";
--X69Y47, nonlinear_LMDPL
constant Tile_X69Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y47, linear_LMDPL
constant Tile_X70Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000010101010011001100110011000000000000000000000000000000001101110111011101";
--X71Y47, linear_LMDPL
constant Tile_X71Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000110011001100110000000000000000";
--X72Y47, nonlinear_LMDPL
constant Tile_X72Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110111000000000000000001100110011001100";
--X73Y47, linear_LMDPL
constant Tile_X73Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100110011001100110000000000000000";
--X74Y47, linear_LMDPL
constant Tile_X74Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000";
--X75Y47, nonlinear_LMDPL
constant Tile_X75Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X76Y47, linear_LMDPL
constant Tile_X76Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X77Y47, linear_LMDPL
constant Tile_X77Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X78Y47, ctrl_to_sec
constant Tile_X78Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y47, combined_WDDL
constant Tile_X79Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y47, combined_WDDL
constant Tile_X80Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y47, ctrl_IO
constant Tile_X81Y47_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y48, W_IO_custom
constant Tile_X0Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y48, linear_LMDPL
constant Tile_X1Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101011010101011111111010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X2Y48, linear_LMDPL
constant Tile_X2Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011";
--X3Y48, nonlinear_LMDPL
constant Tile_X3Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000011001100110011";
--X4Y48, linear_LMDPL
constant Tile_X4Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111111111111110101010010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X5Y48, linear_LMDPL
constant Tile_X5Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010101111111100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001010101010101010";
--X6Y48, nonlinear_LMDPL
constant Tile_X6Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000011001100110011";
--X7Y48, linear_LMDPL
constant Tile_X7Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X8Y48, linear_LMDPL
constant Tile_X8Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X9Y48, nonlinear_LMDPL
constant Tile_X9Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000010101010000000000101010100000000000000001010101010101010010101010101010100000000000000000000000000000000000000000000000000010001000100010000000000000000";
--X10Y48, linear_LMDPL
constant Tile_X10Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X11Y48, linear_LMDPL
constant Tile_X11Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X12Y48, nonlinear_LMDPL
constant Tile_X12Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X13Y48, linear_LMDPL
constant Tile_X13Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000010101010000000000000000010101010000000001111111110101010101010100000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X14Y48, linear_LMDPL
constant Tile_X14Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010101010100000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000100010001000100";
--X15Y48, nonlinear_LMDPL
constant Tile_X15Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X16Y48, linear_LMDPL
constant Tile_X16Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X17Y48, linear_LMDPL
constant Tile_X17Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X18Y48, nonlinear_LMDPL
constant Tile_X18Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111101010101010101000000000000000001010101000000000000000000000000010101010010101010101010100000000101010100001000100010001000000000000000010001000100010000000000000000000";
--X19Y48, linear_LMDPL
constant Tile_X19Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000001111111110101010101010101010101001010101000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X20Y48, linear_LMDPL
constant Tile_X20Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010000000000000000010001000100010000000000010101010000000000000000101110111011101100110011001100110000000000000000";
--X21Y48, nonlinear_LMDPL
constant Tile_X21Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111101010100101010100000000000000001010101000000000000000000000000000000000010001000100010000000000101010100000000000000000100110011001100100000000000000000000000000000000";
--X22Y48, linear_LMDPL
constant Tile_X22Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111011101110111000000000000000000110011001100110";
--X23Y48, linear_LMDPL
constant Tile_X23Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000001010101001010101101010100101010101010101000000000000000000000000111111110000000010101010010101010101010100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X24Y48, nonlinear_LMDPL
constant Tile_X24Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000001010101000000001010101000000000000000000000000001010101010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X25Y48, linear_LMDPL
constant Tile_X25Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111110101010010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X26Y48, linear_LMDPL
constant Tile_X26Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000001010101010101010101010100000000000000000101010101010101000000000000000001100110011001100000000000000000";
--X27Y48, nonlinear_LMDPL
constant Tile_X27Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000001100110011001100110011001100110000000000000000";
--X28Y48, linear_LMDPL
constant Tile_X28Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000001010101101010100000000001010101010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X29Y48, linear_LMDPL
constant Tile_X29Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010101111111100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010110101010000000001011101110111011000000000000000011111111111111110000000000000000";
--X30Y48, nonlinear_LMDPL
constant Tile_X30Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y48, linear_LMDPL
constant Tile_X31Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110100000000000000000000000000000000";
--X32Y48, linear_LMDPL
constant Tile_X32Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101011010101011111111000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000111011101110111001000100010001000000000000000000";
--X33Y48, nonlinear_LMDPL
constant Tile_X33Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101101010100000000000000000000000000000000010101010000000001111111101010101000000000000000000000000010101011010101000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000000000000000000000000000000000000";
--X34Y48, linear_LMDPL
constant Tile_X34Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X35Y48, linear_LMDPL
constant Tile_X35Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000001111111101010101010001000100010000000000000000000000000000000000110111011101110101000100010001000000000000000000";
--X36Y48, nonlinear_LMDPL
constant Tile_X36Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000101010100000000001010101000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X37Y48, linear_LMDPL
constant Tile_X37Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101000000000000000000101010110101010000000000000000000000000000000000000000001010101000000001010101010101010000000000000000000000000000000000101010101010101010101010101010100000000000000001000100010001000000000000000000001110111011101110000000000000000";
--X38Y48, linear_LMDPL
constant Tile_X38Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000010101010010101010101010101010101000000001000100010001000000000000000000000000000000000000000000000000000";
--X39Y48, nonlinear_LMDPL
constant Tile_X39Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y48, linear_LMDPL
constant Tile_X40Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000010101010100010001000100000000000000000000000000000000000000000000000000";
--X41Y48, linear_LMDPL
constant Tile_X41Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010010101010101010100000000101010101101110111011101000000000000000001100110011001100000000000000000";
--X42Y48, nonlinear_LMDPL
constant Tile_X42Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101011010101000000000000000001010101000000000111111110000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X43Y48, linear_LMDPL
constant Tile_X43Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000101010110101010000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000010101011010101010101010000000000000000000000000000000001011101110111011";
--X44Y48, linear_LMDPL
constant Tile_X44Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010000000000000000101010100000000000000000000000000000000001010101000000000000000001010101111111110000000010101010000000000101010100000000101010100000000000000000101010100000000010101010000000000000000000000000000000000000000000000000010101010000000000000000100010001000100000000000000000001011101110111011";
--X45Y48, nonlinear_LMDPL
constant Tile_X45Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X46Y48, linear_LMDPL
constant Tile_X46Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101000000000101010100101010110101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110101000100010001000000000000000000";
--X47Y48, linear_LMDPL
constant Tile_X47Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000010101010000000001111111100000000010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X48Y48, nonlinear_LMDPL
constant Tile_X48Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001011101110111011000000000000000001000100010001000000000000000000";
--X49Y48, linear_LMDPL
constant Tile_X49Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000010101010101010101010101010101010010001000100010000000000000000000000000000000000010101010101010111101110111011100000000000000000";
--X50Y48, linear_LMDPL
constant Tile_X50Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000010101010000000000000000000000000000000000000000111111110000000010101010000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011000100010001000100000000000000000";
--X51Y48, nonlinear_LMDPL
constant Tile_X51Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000101010100000000000000000101010100000000000000001010101000000000101010100000000001010101010001000100010000000000101010100000000000000000100110011001100101000100010001000000000000000000";
--X52Y48, linear_LMDPL
constant Tile_X52Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000011111111101010101010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X53Y48, linear_LMDPL
constant Tile_X53Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001100110011001100";
--X54Y48, nonlinear_LMDPL
constant Tile_X54Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X55Y48, linear_LMDPL
constant Tile_X55Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000110011001100110000000000000000001010101010101010";
--X56Y48, linear_LMDPL
constant Tile_X56Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001111111111111111";
--X57Y48, nonlinear_LMDPL
constant Tile_X57Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111010101000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001011101110111011";
--X58Y48, linear_LMDPL
constant Tile_X58Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000001100110011001100";
--X59Y48, linear_LMDPL
constant Tile_X59Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010010001000100010011111111000000000000000000000000001000100010001000100010001000100000000000000000";
--X60Y48, nonlinear_LMDPL
constant Tile_X60Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101011111111000000000000000001010101000000001010101000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001100110011001100";
--X61Y48, linear_LMDPL
constant Tile_X61Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000010101010010101010101010110101010000000001000100010001000000000000000000000000000000000000000000000000000";
--X62Y48, linear_LMDPL
constant Tile_X62Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000110111011101110100000000000000001010101010101010";
--X63Y48, nonlinear_LMDPL
constant Tile_X63Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X64Y48, linear_LMDPL
constant Tile_X64Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X65Y48, linear_LMDPL
constant Tile_X65Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X66Y48, nonlinear_LMDPL
constant Tile_X66Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y48, linear_LMDPL
constant Tile_X67Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X68Y48, linear_LMDPL
constant Tile_X68Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001000100010001000";
--X69Y48, nonlinear_LMDPL
constant Tile_X69Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001100110011001100";
--X70Y48, linear_LMDPL
constant Tile_X70Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X71Y48, linear_LMDPL
constant Tile_X71Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000011111111000000001010101000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X72Y48, nonlinear_LMDPL
constant Tile_X72Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000100010001000100000000000000000";
--X73Y48, linear_LMDPL
constant Tile_X73Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X74Y48, linear_LMDPL
constant Tile_X74Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000101010100000000000000000010101010000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000110011001100110";
--X75Y48, nonlinear_LMDPL
constant Tile_X75Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001001100110011001";
--X76Y48, linear_LMDPL
constant Tile_X76Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000100010001000100";
--X77Y48, linear_LMDPL
constant Tile_X77Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X78Y48, ctrl_to_sec
constant Tile_X78Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y48, combined_WDDL
constant Tile_X79Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y48, combined_WDDL
constant Tile_X80Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y48, ctrl_IO
constant Tile_X81Y48_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y49, W_IO_custom
constant Tile_X0Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y49, linear_LMDPL
constant Tile_X1Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010111111111010101010101010010101010101010100000000111111110101010101010101000000000000000011101110111011100000000000000000";
--X2Y49, linear_LMDPL
constant Tile_X2Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101011111111100000000010101010101010100000000111111111110111011101110000000000000000000000000000000000000000000000000";
--X3Y49, nonlinear_LMDPL
constant Tile_X3Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000011001100110011";
--X4Y49, linear_LMDPL
constant Tile_X4Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000010101010010001000100010000000000101010100000000000000000110011001100110010001000100010000000000000000000";
--X5Y49, linear_LMDPL
constant Tile_X5Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010101010101010101011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000100010001000100";
--X6Y49, nonlinear_LMDPL
constant Tile_X6Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000011001100110011";
--X7Y49, linear_LMDPL
constant Tile_X7Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000010001000100010000000000000000";
--X8Y49, linear_LMDPL
constant Tile_X8Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000";
--X9Y49, nonlinear_LMDPL
constant Tile_X9Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y49, linear_LMDPL
constant Tile_X10Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111110101010000000001010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X11Y49, linear_LMDPL
constant Tile_X11Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000011111111000000000000000010101010010101010101010100000000000000000111011101110111000000000000000001000100010001000000000000000000";
--X12Y49, nonlinear_LMDPL
constant Tile_X12Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000101010101111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000010001000100010";
--X13Y49, linear_LMDPL
constant Tile_X13Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101010101010000000000000000000000000101010100000000010101010000100010001000100000000101010101011101110111011000000000000000000000000000000001011101110111011";
--X14Y49, linear_LMDPL
constant Tile_X14Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111110101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000101010110101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001101110111011101";
--X15Y49, nonlinear_LMDPL
constant Tile_X15Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000100010001000100";
--X16Y49, linear_LMDPL
constant Tile_X16Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X17Y49, linear_LMDPL
constant Tile_X17Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000100010001000100000000000000000000100010001000100";
--X18Y49, nonlinear_LMDPL
constant Tile_X18Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000111111111010101001010101000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000001100110011001100010001000100010000000000000000";
--X19Y49, linear_LMDPL
constant Tile_X19Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000001010101000000000101010100000000000000000111111110000000010101010101010100000000000000000111111111010101000000000000000000000000010101010010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X20Y49, linear_LMDPL
constant Tile_X20Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101000000001111111100000000000000000000000010101010000000000000000000000000101010101111111100000000000000001010101010101010000000000101010100000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000010001000100010001010101010101010000000000000000";
--X21Y49, nonlinear_LMDPL
constant Tile_X21Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000010001000100010";
--X22Y49, linear_LMDPL
constant Tile_X22Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000001010101001010101010001000100010010101010000000000000000000000000101010101010101001000100010001000000000000000000";
--X23Y49, linear_LMDPL
constant Tile_X23Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000101010100000000000000000000000000000000010101010000000001010101001010101101010100000000000000000000000001010101010101010101010100000000010101010000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000101110111011101100000000000000001101110111011101";
--X24Y49, nonlinear_LMDPL
constant Tile_X24Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000010101010010001000100010000000000101010100000000000000000000000000000000001100110011001100000000000000000";
--X25Y49, linear_LMDPL
constant Tile_X25Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000001010101000000000000000000000000010101010000000000000000000000000010101011010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X26Y49, linear_LMDPL
constant Tile_X26Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101011111111110101010010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X27Y49, nonlinear_LMDPL
constant Tile_X27Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X28Y49, linear_LMDPL
constant Tile_X28Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000101010101111111100000000000100010001000111111111000000001000100010001000000000000000000000000000000000000100010001000100";
--X29Y49, linear_LMDPL
constant Tile_X29Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001110111011101110";
--X30Y49, nonlinear_LMDPL
constant Tile_X30Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X31Y49, linear_LMDPL
constant Tile_X31Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000001010101010101010101010100000000000000000000000000000000000000000000000000110011001100110000000000000000";
--X32Y49, linear_LMDPL
constant Tile_X32Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000101010101111111101010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000110011001100110000000000000000010001000100010000000000000000000";
--X33Y49, nonlinear_LMDPL
constant Tile_X33Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X34Y49, linear_LMDPL
constant Tile_X34Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000001010101000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000001000100010001000100010001000100000000000000000";
--X35Y49, linear_LMDPL
constant Tile_X35Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X36Y49, nonlinear_LMDPL
constant Tile_X36Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000001010101000000000000000000000000010101010000100010001000100000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X37Y49, linear_LMDPL
constant Tile_X37Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111010101010101010000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X38Y49, linear_LMDPL
constant Tile_X38Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000001010101010101010101010101111111110101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X39Y49, nonlinear_LMDPL
constant Tile_X39Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X40Y49, linear_LMDPL
constant Tile_X40Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000011111111010101010101010100000000101010101100110011001100000000000000000011011101110111010000000000000000";
--X41Y49, linear_LMDPL
constant Tile_X41Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000001010101000000000000000000000000000000000010001000100010000000000111111110000000000000000001000100010001010111011101110110000000000000000";
--X42Y49, nonlinear_LMDPL
constant Tile_X42Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101011111111000000000000000000000000000000000000000010101010000100010001000100000000010101010010001000100010000000000000000000000000000000000101010101010101";
--X43Y49, linear_LMDPL
constant Tile_X43Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000101010110101010000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000001100110011001100000000000000000000000000000000";
--X44Y49, linear_LMDPL
constant Tile_X44Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000010101010010101010000000000000000101010100000000000000000101010100000000010101010010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X45Y49, nonlinear_LMDPL
constant Tile_X45Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000100110011001100100000000000000001010101010101010";
--X46Y49, linear_LMDPL
constant Tile_X46Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000111111110101010100000000010101011010101010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101110111011101100000000000000001000100010001000";
--X47Y49, linear_LMDPL
constant Tile_X47Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110010111011101110110000000000000000";
--X48Y49, nonlinear_LMDPL
constant Tile_X48Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X49Y49, linear_LMDPL
constant Tile_X49Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010000000000000000010101010101010101010101010101010000000000000000000000000000000000000000000000000011001100110011000000000000000000010001000100010";
--X50Y49, linear_LMDPL
constant Tile_X50Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X51Y49, nonlinear_LMDPL
constant Tile_X51Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001010101000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000000000000000000000000010101010000000000000000101110111011101100000000000000001100110011001100";
--X52Y49, linear_LMDPL
constant Tile_X52Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X53Y49, linear_LMDPL
constant Tile_X53Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X54Y49, nonlinear_LMDPL
constant Tile_X54Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X55Y49, linear_LMDPL
constant Tile_X55Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010101010100101010111111111000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X56Y49, linear_LMDPL
constant Tile_X56Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X57Y49, nonlinear_LMDPL
constant Tile_X57Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001000100010001000";
--X58Y49, linear_LMDPL
constant Tile_X58Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101010101010000000000000000001010101000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000100010001000100000000000000000001110111011101110";
--X59Y49, linear_LMDPL
constant Tile_X59Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010010001000100010010101010101010100000000000000000100010001000100000110011001100110000000000000000";
--X60Y49, nonlinear_LMDPL
constant Tile_X60Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y49, linear_LMDPL
constant Tile_X61Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000101010110101010000000000000000000000000000000000000000000000000101010100000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001010101010101010";
--X62Y49, linear_LMDPL
constant Tile_X62Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000000000000010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X63Y49, nonlinear_LMDPL
constant Tile_X63Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101110111011101100000000000000001001100110011001";
--X64Y49, linear_LMDPL
constant Tile_X64Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X65Y49, linear_LMDPL
constant Tile_X65Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000101010100000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111011101110";
--X66Y49, nonlinear_LMDPL
constant Tile_X66Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000111111110000000000000000010001000100010000000000000000000000000000000000101110111011101110001000100010000000000000000000";
--X67Y49, linear_LMDPL
constant Tile_X67Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X68Y49, linear_LMDPL
constant Tile_X68Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010101010101010110101010000000001100110011001100000000000000000010101010101010100000000000000000";
--X69Y49, nonlinear_LMDPL
constant Tile_X69Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X70Y49, linear_LMDPL
constant Tile_X70Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000010101010101010101010101000000000010101010000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001001000100010001000000000000000000";
--X71Y49, linear_LMDPL
constant Tile_X71Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000111111110000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X72Y49, nonlinear_LMDPL
constant Tile_X72Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001000100010001000";
--X73Y49, linear_LMDPL
constant Tile_X73Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000010001000100010";
--X74Y49, linear_LMDPL
constant Tile_X74Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000001000100010001";
--X75Y49, nonlinear_LMDPL
constant Tile_X75Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X76Y49, linear_LMDPL
constant Tile_X76Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X77Y49, linear_LMDPL
constant Tile_X77Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000111111111000000000111011101110111000000000000000000000000000000000000000000000000";
--X78Y49, ctrl_to_sec
constant Tile_X78Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y49, combined_WDDL
constant Tile_X79Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y49, combined_WDDL
constant Tile_X80Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y49, ctrl_IO
constant Tile_X81Y49_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y50, W_IO_custom
constant Tile_X0Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y50, linear_LMDPL
constant Tile_X1Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101011111111000000000000000000000000101010101010101010101010010001000100010000000000000000000000000000000000010001000100010000100010001000100000000000000000";
--X2Y50, linear_LMDPL
constant Tile_X2Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000010101010101010100000000000000000010101010101010100000000000000001101110111011101000000000000000010111011101110110000000000000000";
--X3Y50, nonlinear_LMDPL
constant Tile_X3Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000010001000100010";
--X4Y50, linear_LMDPL
constant Tile_X4Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010101010101010100000000000000001000100010001000000000000000000010011001100110010000000000000000";
--X5Y50, linear_LMDPL
constant Tile_X5Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010111111111010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001001100110011001";
--X6Y50, nonlinear_LMDPL
constant Tile_X6Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X7Y50, linear_LMDPL
constant Tile_X7Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000111011101110111";
--X8Y50, linear_LMDPL
constant Tile_X8Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101011111111000000000000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X9Y50, nonlinear_LMDPL
constant Tile_X9Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000101010100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001001100110011001000000000000000000000000000000001100110011001100";
--X10Y50, linear_LMDPL
constant Tile_X10Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000111111111010101010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X11Y50, linear_LMDPL
constant Tile_X11Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000011101110111011100000000000000001100110011001100";
--X12Y50, nonlinear_LMDPL
constant Tile_X12Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000011111111000000000101010100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000111011101110111";
--X13Y50, linear_LMDPL
constant Tile_X13Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111111111111000000001010101010101010000000001010101010101010101010100000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000001101110111011101";
--X14Y50, linear_LMDPL
constant Tile_X14Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010101010100000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X15Y50, nonlinear_LMDPL
constant Tile_X15Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000001010101000000000000000000101010100000000000000000000000001010101101010100000000000000000010101010101010100000000000000000000000000000000000000000000000000010001000100010000000000000000";
--X16Y50, linear_LMDPL
constant Tile_X16Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000001010101000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X17Y50, linear_LMDPL
constant Tile_X17Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000000000000000000000110011001100110000000000000000";
--X18Y50, nonlinear_LMDPL
constant Tile_X18Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000001010101000000000101010100101010100000000000000001010101000000000111111110000000010101010010001000100010000000000101010100000000000000000000100010001000110001000100010000000000000000000";
--X19Y50, linear_LMDPL
constant Tile_X19Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010110101010111111110101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000001110111011101110000000000000000";
--X20Y50, linear_LMDPL
constant Tile_X20Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000000000000000010101010101010101010101000000000000000000000000000000000101010100101010101010101000100010001000100000000000000000110011001100110000000000000000000000000000000001100110011001100";
--X21Y50, nonlinear_LMDPL
constant Tile_X21Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101000000000000000000000000001010101111111111010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000000001000100010001";
--X22Y50, linear_LMDPL
constant Tile_X22Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101000000000000000000101010100000000000000001111111100000000000000000101010110101010010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X23Y50, linear_LMDPL
constant Tile_X23Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000001010101010101010101010100000000010101010000000000000000000000000101010100000000010101010010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X24Y50, nonlinear_LMDPL
constant Tile_X24Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000001010101000000000101010100000000001010101010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X25Y50, linear_LMDPL
constant Tile_X25Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000011111111000000001010101000000000101010101010101010101010010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X26Y50, linear_LMDPL
constant Tile_X26Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111111111111010101010101010010101010101010110101010000000000100010001000100000000000000000011001100110011000000000000000000";
--X27Y50, nonlinear_LMDPL
constant Tile_X27Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000110011001100110";
--X28Y50, linear_LMDPL
constant Tile_X28Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010101010101010101010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X29Y50, linear_LMDPL
constant Tile_X29Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111111110101010100000000010001000100010000000000000000000000000000000000110011001100110011111111111111110000000000000000";
--X30Y50, nonlinear_LMDPL
constant Tile_X30Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X31Y50, linear_LMDPL
constant Tile_X31Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010010101011111111100000000101010100000000000000000000000001010101000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000101110111011101111001100110011000000000000000000";
--X32Y50, linear_LMDPL
constant Tile_X32Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000000000000011111111010101010101010100000000000000001010101010101010000000000000000001110111011101110000000000000000";
--X33Y50, nonlinear_LMDPL
constant Tile_X33Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100101010111111111000000001010101000000000000000000000000000000000010101010101010100000000101010100011001100110011000000000000000001000100010001000000000000000000";
--X34Y50, linear_LMDPL
constant Tile_X34Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X35Y50, linear_LMDPL
constant Tile_X35Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001111111100000000010101010000000000000000111111110000000010101010000000000000000000000000101010100000000000000000000100010001000101010101000000000000000000000000000000000000000000000000000000001000100010001000";
--X36Y50, nonlinear_LMDPL
constant Tile_X36Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000010101010000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001010101010101010";
--X37Y50, linear_LMDPL
constant Tile_X37Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001111111101010101010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111111010101010101010010001000100010000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X38Y50, linear_LMDPL
constant Tile_X38Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000010101010000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101010101010010101010101010100000000010101010000000000000000000000000000000011111111111111110000000000000000";
--X39Y50, nonlinear_LMDPL
constant Tile_X39Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000011111111101010100000000000000000111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010101010000000010101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X40Y50, linear_LMDPL
constant Tile_X40Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X41Y50, linear_LMDPL
constant Tile_X41Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000010101010000100010001000100000000101010100011001100110011000000000000000000000000000000000110011001100110";
--X42Y50, nonlinear_LMDPL
constant Tile_X42Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000001010101010101010000000000000000010101010000000000000000000000000010101010000000000000000101010101010101000000000000000000000000000000000";
--X43Y50, linear_LMDPL
constant Tile_X43Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000011111111111111110000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000101010100000000010101010000000000000000000000000101010100000000000000000011001100110011000000000000000000000000000000000";
--X44Y50, linear_LMDPL
constant Tile_X44Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000101010100000000000000000000000010101010000000000101010110101010010001000100010000000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X45Y50, nonlinear_LMDPL
constant Tile_X45Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X46Y50, linear_LMDPL
constant Tile_X46Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111111010101010101010000000000000000000000000101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001101110111011101";
--X47Y50, linear_LMDPL
constant Tile_X47Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001010101010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000101010101010101";
--X48Y50, nonlinear_LMDPL
constant Tile_X48Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101001010101000000000000000000000000101010100000000010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X49Y50, linear_LMDPL
constant Tile_X49Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010101010101000000000010101010101010110101010111111111010101010101010000000000000000011011101110111010000000000000000";
--X50Y50, linear_LMDPL
constant Tile_X50Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000010101011010101010101010010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X51Y50, nonlinear_LMDPL
constant Tile_X51Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000001010101001010101000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010101010100000000000000000000100010001000100000000101010101101110111011101000000000000000000000000000000000100010001000100";
--X52Y50, linear_LMDPL
constant Tile_X52Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010101111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100101010110101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000011101110111011111011101110111010000000000000000";
--X53Y50, linear_LMDPL
constant Tile_X53Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010111111111000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X54Y50, nonlinear_LMDPL
constant Tile_X54Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X55Y50, linear_LMDPL
constant Tile_X55Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101010101010101010100101010100000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000";
--X56Y50, linear_LMDPL
constant Tile_X56Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X57Y50, nonlinear_LMDPL
constant Tile_X57Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X58Y50, linear_LMDPL
constant Tile_X58Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X59Y50, linear_LMDPL
constant Tile_X59Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010010101010101010100000000000000000011001100110011000000000000000001010101010101010000000000000000";
--X60Y50, nonlinear_LMDPL
constant Tile_X60Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000100010001000100";
--X61Y50, linear_LMDPL
constant Tile_X61Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000000000000000000011111111101010100000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001101110111011101";
--X62Y50, linear_LMDPL
constant Tile_X62Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010101010101000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010101010101010101000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X63Y50, nonlinear_LMDPL
constant Tile_X63Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000011001100110011";
--X64Y50, linear_LMDPL
constant Tile_X64Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X65Y50, linear_LMDPL
constant Tile_X65Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000000100010001000101000100010001000000000000000000";
--X66Y50, nonlinear_LMDPL
constant Tile_X66Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000001000100010001";
--X67Y50, linear_LMDPL
constant Tile_X67Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000011001100110011";
--X68Y50, linear_LMDPL
constant Tile_X68Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000100010001000110101010000000000100010001000100000000000000000000000000000000001011101110111011";
--X69Y50, nonlinear_LMDPL
constant Tile_X69Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000010101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001011101110111011";
--X70Y50, linear_LMDPL
constant Tile_X70Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X71Y50, linear_LMDPL
constant Tile_X71Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000101010101010101000000000000000000000000010101010010101010000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X72Y50, nonlinear_LMDPL
constant Tile_X72Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X73Y50, linear_LMDPL
constant Tile_X73Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001100110011001100";
--X74Y50, linear_LMDPL
constant Tile_X74Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000111111110000000000000000000000001010101010101010010101010000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000110011001100110000000000000000";
--X75Y50, nonlinear_LMDPL
constant Tile_X75Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000111111110101010110101010101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X76Y50, linear_LMDPL
constant Tile_X76Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000001000100010001000000000000000001100110011001100";
--X77Y50, linear_LMDPL
constant Tile_X77Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000111011101110111";
--X78Y50, ctrl_to_sec
constant Tile_X78Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y50, combined_WDDL
constant Tile_X79Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y50, combined_WDDL
constant Tile_X80Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y50, ctrl_IO
constant Tile_X81Y50_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y51, W_IO_custom
constant Tile_X0Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y51, linear_LMDPL
constant Tile_X1Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010010101010101010100000000000000001110111011101110000000000000000010001000100010000000000000000000";
--X2Y51, linear_LMDPL
constant Tile_X2Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000010101010101010100000000000000000010001000100010000000000111111110000000000000000000100010001000111101110111011100000000000000000";
--X3Y51, nonlinear_LMDPL
constant Tile_X3Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000100010001000100000000000000000001000100010001000000000000000000000000000000000101010101010101";
--X4Y51, linear_LMDPL
constant Tile_X4Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101111111100000000010001000100010000000000000000000000000000000000011001100110011011101110111011100000000000000000";
--X5Y51, linear_LMDPL
constant Tile_X5Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010101010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X6Y51, nonlinear_LMDPL
constant Tile_X6Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000011001100110011";
--X7Y51, linear_LMDPL
constant Tile_X7Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X8Y51, linear_LMDPL
constant Tile_X8Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X9Y51, nonlinear_LMDPL
constant Tile_X9Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000010101010000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000000010001000100010000000000000000";
--X10Y51, linear_LMDPL
constant Tile_X10Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000001010101010101010010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X11Y51, linear_LMDPL
constant Tile_X11Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X12Y51, nonlinear_LMDPL
constant Tile_X12Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000001111111110101010010001000100010000000000000000000000000000000000100110011001100100100010001000100000000000000000";
--X13Y51, linear_LMDPL
constant Tile_X13Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010101111111101010101000100010001000100000000101010101010101010101010000000000000000000000000000000000000000000000000";
--X14Y51, linear_LMDPL
constant Tile_X14Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000001010101000000000000000000000000101010100000000000000000010101010101010100000000101010101000100010001000000000000000000001000100010001000000000000000000";
--X15Y51, nonlinear_LMDPL
constant Tile_X15Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001011101110111011";
--X16Y51, linear_LMDPL
constant Tile_X16Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000110011001100110";
--X17Y51, linear_LMDPL
constant Tile_X17Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000000110011001100110000000000000000";
--X18Y51, nonlinear_LMDPL
constant Tile_X18Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000111111110000000010101010000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000100010001000100011001100110011000000000000000000";
--X19Y51, linear_LMDPL
constant Tile_X19Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101010101010000000000101010100000000000000001010101000000000000000000101010100000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X20Y51, linear_LMDPL
constant Tile_X20Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000010101010000000000000000000000000101010110101010101010100101010100000000000000000000000000000000111111111010101010101010010101010101010100000000000000000101010101010101000000000000000001100110011001100000000000000000";
--X21Y51, nonlinear_LMDPL
constant Tile_X21Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000001111111100000000101010100000000010101010000000001010101000000000000000000000000000000000010001000100010000000000101010100000000000000000101110111011101101110111011101110000000000000000";
--X22Y51, linear_LMDPL
constant Tile_X22Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100101010100000000000000001010101011111111000000000000000000000000000000000000000011111111000000001010101000000000101010100101010100000000101010100000000000000000000000001010101010101010010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X23Y51, linear_LMDPL
constant Tile_X23Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010101010101010101010101010100000000010101010000000000000000000000000111111110000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X24Y51, nonlinear_LMDPL
constant Tile_X24Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000001010101010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000001010101010001000100010000000000101010100000000000000000110011001100110000000000000000000000000000000000";
--X25Y51, linear_LMDPL
constant Tile_X25Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010101010101000000000010101011010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000010101011010101010101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X26Y51, linear_LMDPL
constant Tile_X26Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101011111111010001000100010000000000111111110000000000000000010001000100010000000000000000000000000000000000";
--X27Y51, nonlinear_LMDPL
constant Tile_X27Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000011001100110011";
--X28Y51, linear_LMDPL
constant Tile_X28Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000011111111010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X29Y51, linear_LMDPL
constant Tile_X29Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000001010101000100010001000110101010000000000000000000000000000000000000000000000000000000001000100010001000";
--X30Y51, nonlinear_LMDPL
constant Tile_X30Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101010101010100000000000000001001100110011001000000000000000000110011001100110000000000000000";
--X31Y51, linear_LMDPL
constant Tile_X31Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101010101010101010100000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000101010101010101010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X32Y51, linear_LMDPL
constant Tile_X32Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000100010001000101010101000000000000000000000000000000000000000000000000000000001000100010001000";
--X33Y51, nonlinear_LMDPL
constant Tile_X33Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000111111110000000001010101000000000000000000000000000000001010101000000000101010101010101000000000000000001010101000000000010101010000000000000000010001000100010000000000000000000000000000000000101110111011101100100010001000100000000000000000";
--X34Y51, linear_LMDPL
constant Tile_X34Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000101010100000000111111110000000000000000000000000000000010101010000000000101010110101010000000000000000000000000000000000000000001010101010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X35Y51, linear_LMDPL
constant Tile_X35Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100101010100000000010101010101010100000000000000000000000000000000000000000000000010101010101010100000000000000000";
--X36Y51, nonlinear_LMDPL
constant Tile_X36Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000010101010000000001010101000000000010101010101010110101010010001000100010000000000101010100000000000000000110011001100110010001000100010000000000000000000";
--X37Y51, linear_LMDPL
constant Tile_X37Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000001010101000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000111111111010101010101010010101010101010101010101111111111100110011001100000000000000000010001000100010000000000000000000";
--X38Y51, linear_LMDPL
constant Tile_X38Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000101010100000000001010101000000001010101000000000000000001111111100000000000000000000000000000000000000001010101010101010101010101111111110101010010101010101010100000000000000001111111111111111000000000000000000110011001100110000000000000000";
--X39Y51, nonlinear_LMDPL
constant Tile_X39Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000001010101000000000000000000000000010101010000100010001000100000000010101011100110011001100000000000000000000000000000000001000100010001000";
--X40Y51, linear_LMDPL
constant Tile_X40Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111101010100000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010010101010101010100000000101010100010001000100010000000000000000010111011101110110000000000000000";
--X41Y51, linear_LMDPL
constant Tile_X41Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000111111111010101010101010000000001010101001010101000000000000000010101010000000000000000000000000101010100000000000000000101010101010101000000000000000000010001000100010";
--X42Y51, nonlinear_LMDPL
constant Tile_X42Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010101010101000000000000000000110011001100110";
--X43Y51, linear_LMDPL
constant Tile_X43Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010101010100000000010101010000000000000000010101010111111110101010110101010000000000000000000000000101010100000000010101010000000000000000000000000010101010000000000000000110011001100110000000000000000001010101010101010";
--X44Y51, linear_LMDPL
constant Tile_X44Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000011111111000000000101010100000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101010111011101110110000000000000000";
--X45Y51, nonlinear_LMDPL
constant Tile_X45Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000001010101000000000000000000000000010101010000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X46Y51, linear_LMDPL
constant Tile_X46Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101011111111101010101010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X47Y51, linear_LMDPL
constant Tile_X47Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X48Y51, nonlinear_LMDPL
constant Tile_X48Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X49Y51, linear_LMDPL
constant Tile_X49Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101010101000000000010101010101010100000000000000001000100010001000000000000000000011011101110111010000000000000000";
--X50Y51, linear_LMDPL
constant Tile_X50Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010101010101000000000000100010001000111111111000000001010101010101010000000000000000000000000000000000011001100110011";
--X51Y51, nonlinear_LMDPL
constant Tile_X51Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000000100010001000100";
--X52Y51, linear_LMDPL
constant Tile_X52Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X53Y51, linear_LMDPL
constant Tile_X53Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000000000001010101000000000101010101010101000000000010001000100010000000000000000000000000000000000101110111011101110001000100010000000000000000000";
--X54Y51, nonlinear_LMDPL
constant Tile_X54Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000110011001100110";
--X55Y51, linear_LMDPL
constant Tile_X55Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000010101010000000000000000111111111010101000000000000000001010101001010101101010100000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X56Y51, linear_LMDPL
constant Tile_X56Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X57Y51, nonlinear_LMDPL
constant Tile_X57Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X58Y51, linear_LMDPL
constant Tile_X58Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000000000000000000000000000000000000111111111111111100000000000000001011101110111011";
--X59Y51, linear_LMDPL
constant Tile_X59Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000101010101010101010101010010101010101010110101010101010101101110111011101000000000000000000100010001000100000000000000000";
--X60Y51, nonlinear_LMDPL
constant Tile_X60Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000001001100110011001";
--X61Y51, linear_LMDPL
constant Tile_X61Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000010101010000000000000000010101010000000000000000000000000100110011001100100000000000000000010001000100010";
--X62Y51, linear_LMDPL
constant Tile_X62Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000111011101110111000000000000000000000000000000000";
--X63Y51, nonlinear_LMDPL
constant Tile_X63Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X64Y51, linear_LMDPL
constant Tile_X64Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X65Y51, linear_LMDPL
constant Tile_X65Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000";
--X66Y51, nonlinear_LMDPL
constant Tile_X66Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X67Y51, linear_LMDPL
constant Tile_X67Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X68Y51, linear_LMDPL
constant Tile_X68Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X69Y51, nonlinear_LMDPL
constant Tile_X69Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X70Y51, linear_LMDPL
constant Tile_X70Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X71Y51, linear_LMDPL
constant Tile_X71Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000101010100000000000000000000000001010101000000000010101011010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100000000000000000000100010001000100000000000000000";
--X72Y51, nonlinear_LMDPL
constant Tile_X72Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010111111110000000000000000000000001010101000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X73Y51, linear_LMDPL
constant Tile_X73Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101000000001111111110101010000000000000000000000000000000000101010111111111101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000110011001100110000000000000000000000000000000000";
--X74Y51, linear_LMDPL
constant Tile_X74Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X75Y51, nonlinear_LMDPL
constant Tile_X75Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010";
--X76Y51, linear_LMDPL
constant Tile_X76Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111011101110111000000000000000001000100010001000";
--X77Y51, linear_LMDPL
constant Tile_X77Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001011101110111011";
--X78Y51, ctrl_to_sec
constant Tile_X78Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y51, combined_WDDL
constant Tile_X79Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y51, combined_WDDL
constant Tile_X80Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y51, ctrl_IO
constant Tile_X81Y51_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y52, W_IO_custom
constant Tile_X0Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000";
--X1Y52, linear_LMDPL
constant Tile_X1Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111111010101010101010000000000000000011111111000000000000000000000000010101010101010100000000000000000001000100010001";
--X2Y52, linear_LMDPL
constant Tile_X2Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000010111011101110110000000000000000";
--X3Y52, nonlinear_LMDPL
constant Tile_X3Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X4Y52, linear_LMDPL
constant Tile_X4Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X5Y52, linear_LMDPL
constant Tile_X5Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001101110111011101";
--X6Y52, nonlinear_LMDPL
constant Tile_X6Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000101010101010101";
--X7Y52, linear_LMDPL
constant Tile_X7Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X8Y52, linear_LMDPL
constant Tile_X8Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001111111111111111";
--X9Y52, nonlinear_LMDPL
constant Tile_X9Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y52, linear_LMDPL
constant Tile_X10Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X11Y52, linear_LMDPL
constant Tile_X11Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X12Y52, nonlinear_LMDPL
constant Tile_X12Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110010111011101110110000000000000000";
--X13Y52, linear_LMDPL
constant Tile_X13Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101010101010000000001010101010101010101010100000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X14Y52, linear_LMDPL
constant Tile_X14Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010101010101010101000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X15Y52, nonlinear_LMDPL
constant Tile_X15Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001111111101010101101010101010101001010101000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000101110111011101110001000100010000000000000000000";
--X16Y52, linear_LMDPL
constant Tile_X16Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001000100010001000000000000000000001110111011101110000000000000000";
--X17Y52, linear_LMDPL
constant Tile_X17Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000010101010010101010101010110101010000000000000000000000000000000000000000001100110011001100000000000000000";
--X18Y52, nonlinear_LMDPL
constant Tile_X18Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000010101011010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000101010100000000000000001010101000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000000000000000000000001000100010001";
--X19Y52, linear_LMDPL
constant Tile_X19Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100000000010101010010101011111111111111111000000000000000010101010000000000101010101010101000000000000000000000000000000000000000000000000010101010101010100000000101010100011001100110011000000000000000000100010001000100000000000000000";
--X20Y52, linear_LMDPL
constant Tile_X20Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010101010101010101011111111000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X21Y52, nonlinear_LMDPL
constant Tile_X21Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000010101010000000000000000111111110000000000000000000000000000000001010101101010100000000000000000000000000000000010101010010101010000000010101010000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000001100110011001100";
--X22Y52, linear_LMDPL
constant Tile_X22Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111101010101111111100000000000000000000000000000000000000000101010100000000101010100000000000000000000000001010101000000000010101010101010100000000000000000000000000000000000000001010101010101010000100010001000110101010000000000100010001000100000000000000000000000000000000001111111111111111";
--X23Y52, linear_LMDPL
constant Tile_X23Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X24Y52, nonlinear_LMDPL
constant Tile_X24Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010110101010101010100000000000000000000000001010101000000000000000000000000000000000000000001010101000000000101010100101010101010101010001000100010000000000000000000000000000000000101110111011101110101010101010100000000000000000";
--X25Y52, linear_LMDPL
constant Tile_X25Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000101010100101010110101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X26Y52, linear_LMDPL
constant Tile_X26Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000011111111101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000001010101010101010101010100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X27Y52, nonlinear_LMDPL
constant Tile_X27Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101011010101000000000000000000000000011111111000000001010101000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000100010001000100000000000000001100110011001100000000000000000000000000000000000110011001100110";
--X28Y52, linear_LMDPL
constant Tile_X28Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101011010101011111111000100010001000110101010000000001010101010101010000000000000000000000000000000000000000000000000";
--X29Y52, linear_LMDPL
constant Tile_X29Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001111111110101010010101010101010100000000000000000110011001100110000000000000000000110011001100110000000000000000";
--X30Y52, nonlinear_LMDPL
constant Tile_X30Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101000100010001000100000000000000000";
--X31Y52, linear_LMDPL
constant Tile_X31Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010101010100000000000000000101010100000000011111111000000001010101000000000000000000000000000000000010101011010101010101010010001000100010000000000000000000000000000000000101010101010101000000000000000000000000000000000";
--X32Y52, linear_LMDPL
constant Tile_X32Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000111011101110111010101010101010100000000000000000";
--X33Y52, nonlinear_LMDPL
constant Tile_X33Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000010101010000000000000000001010101000000000000000011111111000000001010101000000000101010100000000000000000000000001010101000000000010101010000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000000010001000100010";
--X34Y52, linear_LMDPL
constant Tile_X34Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000101010100101010110101010000000000000000000000000111111110101010100000000010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X35Y52, linear_LMDPL
constant Tile_X35Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111101010100101010101010101010101010000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001101110111011101";
--X36Y52, nonlinear_LMDPL
constant Tile_X36Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000010101010000000001010101000000000101010101010101001010101010001000100010000000000010101010000000000000000110011001100110000000000000000000000000000000000";
--X37Y52, linear_LMDPL
constant Tile_X37Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010101010101111111100000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010101010101000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001111111111111111";
--X38Y52, linear_LMDPL
constant Tile_X38Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000101010101010101010101010000000000000000011001100110011000000000000000000";
--X39Y52, nonlinear_LMDPL
constant Tile_X39Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000101010100000000010101010000100010001000100000000010101011000100010001000000000000000000000000000000000000000000000000000";
--X40Y52, linear_LMDPL
constant Tile_X40Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000010101010101010100000000111111110000000000000000000000000000000000100010001000100000000000000000";
--X41Y52, linear_LMDPL
constant Tile_X41Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000100010001000100000000010101010011001100110011000000000000000000000000000000001100110011001100";
--X42Y52, nonlinear_LMDPL
constant Tile_X42Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100101010110101010000000001010101010101010000000000000000010101010010001000100010000000000101010100000000000000000110111011101110111001100110011000000000000000000";
--X43Y52, linear_LMDPL
constant Tile_X43Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000010101010000000000000000000000000000000010101010101010100000000010101010000000001010101010101010101010100101010110101010000000000000000000000000101010101010101010101010000100010001000100000000000000001011101110111011000000000000000000000000000000001000100010001000";
--X44Y52, linear_LMDPL
constant Tile_X44Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000111111110000000010101010000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X45Y52, nonlinear_LMDPL
constant Tile_X45Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101011111111101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000110011001100110";
--X46Y52, linear_LMDPL
constant Tile_X46Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111111010101000000000010101011010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X47Y52, linear_LMDPL
constant Tile_X47Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000001011101110111011";
--X48Y52, nonlinear_LMDPL
constant Tile_X48Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X49Y52, linear_LMDPL
constant Tile_X49Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000010001000100010000000000101010100000000000000000010101010101010110111011101110110000000000000000";
--X50Y52, linear_LMDPL
constant Tile_X50Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010110101010000000001010101000000000101010101010101000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X51Y52, nonlinear_LMDPL
constant Tile_X51Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101010101010111111110000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000000100010001000100";
--X52Y52, linear_LMDPL
constant Tile_X52Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X53Y52, linear_LMDPL
constant Tile_X53Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101001010101101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X54Y52, nonlinear_LMDPL
constant Tile_X54Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000";
--X55Y52, linear_LMDPL
constant Tile_X55Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101";
--X56Y52, linear_LMDPL
constant Tile_X56Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X57Y52, nonlinear_LMDPL
constant Tile_X57Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X58Y52, linear_LMDPL
constant Tile_X58Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101011111111000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000101110111011101100000000000000000011001100110011";
--X59Y52, linear_LMDPL
constant Tile_X59Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000100010001000100000000000000001111111111111111000000000000000000000000000000000010001000100010";
--X60Y52, nonlinear_LMDPL
constant Tile_X60Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000010101010111111110000000000000000000000001010101001010101000000000000000000000000000000001010101000000000000000000000000001010101000000000000000000000000000000000000000000000000110011001100110000000000000000001010101010101010";
--X61Y52, linear_LMDPL
constant Tile_X61Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101010101010000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000001010101010101010";
--X62Y52, linear_LMDPL
constant Tile_X62Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101011111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011000000000000000001010101010101010";
--X63Y52, nonlinear_LMDPL
constant Tile_X63Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000001010101010101010";
--X64Y52, linear_LMDPL
constant Tile_X64Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000101010100000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X65Y52, linear_LMDPL
constant Tile_X65Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100";
--X66Y52, nonlinear_LMDPL
constant Tile_X66Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000001000100010001000";
--X67Y52, linear_LMDPL
constant Tile_X67Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X68Y52, linear_LMDPL
constant Tile_X68Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000010101010010001000100010010101010000000000000000000000000101010101010101000010001000100010000000000000000";
--X69Y52, nonlinear_LMDPL
constant Tile_X69Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X70Y52, linear_LMDPL
constant Tile_X70Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001110111011101110";
--X71Y52, linear_LMDPL
constant Tile_X71Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X72Y52, nonlinear_LMDPL
constant Tile_X72Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X73Y52, linear_LMDPL
constant Tile_X73Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000010101010101010100000000000000000000000001010101000000000111111110000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X74Y52, linear_LMDPL
constant Tile_X74Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X75Y52, nonlinear_LMDPL
constant Tile_X75Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X76Y52, linear_LMDPL
constant Tile_X76Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000011001100110011";
--X77Y52, linear_LMDPL
constant Tile_X77Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001111111111111111000000000000000000000000000000000001000100010001";
--X78Y52, ctrl_to_sec
constant Tile_X78Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y52, combined_WDDL
constant Tile_X79Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y52, combined_WDDL
constant Tile_X80Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y52, ctrl_IO
constant Tile_X81Y52_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y53, W_IO_custom
constant Tile_X0Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000";
--X1Y53, linear_LMDPL
constant Tile_X1Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000010101010010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X2Y53, linear_LMDPL
constant Tile_X2Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000000000000000010101010000000001010101000000000010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X3Y53, nonlinear_LMDPL
constant Tile_X3Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X4Y53, linear_LMDPL
constant Tile_X4Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101011111111000000000000000000000000000000001010101000000000010101010101010100000000000000001101110111011101000000000000000011001100110011000000000000000000";
--X5Y53, linear_LMDPL
constant Tile_X5Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000001010101010101010";
--X6Y53, nonlinear_LMDPL
constant Tile_X6Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000110011001100110";
--X7Y53, linear_LMDPL
constant Tile_X7Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000110011001100110000000000000000000010001000100010";
--X8Y53, linear_LMDPL
constant Tile_X8Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000001000100010001";
--X9Y53, nonlinear_LMDPL
constant Tile_X9Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y53, linear_LMDPL
constant Tile_X10Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111111010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X11Y53, linear_LMDPL
constant Tile_X11Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000001100110011001100000000000000000011011101110111010000000000000000";
--X12Y53, nonlinear_LMDPL
constant Tile_X12Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000010101011111111100000000101010100000000000000000000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000001100110011001100010001000100010000000000000000";
--X13Y53, linear_LMDPL
constant Tile_X13Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110111011101110111001100110011000000000000000000";
--X14Y53, linear_LMDPL
constant Tile_X14Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000001010101010101010";
--X15Y53, nonlinear_LMDPL
constant Tile_X15Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101011111111101010101010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010011001100110010000000000000000";
--X16Y53, linear_LMDPL
constant Tile_X16Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000100010001000111111111000000000011001100110011000000000000000000000000000000000011001100110011";
--X17Y53, linear_LMDPL
constant Tile_X17Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X18Y53, nonlinear_LMDPL
constant Tile_X18Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000001010101001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X19Y53, linear_LMDPL
constant Tile_X19Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010000000000000000001010101000000001010101000000000000000001111111100000000010101010101010100000000000000000000000000000000000000000000000001110111011101110000000000000000";
--X20Y53, linear_LMDPL
constant Tile_X20Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001000100010001000000000000000000001010101010101010000000000000000";
--X21Y53, nonlinear_LMDPL
constant Tile_X21Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001111111110101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000100110011001100100000000000000000000000000000000";
--X22Y53, linear_LMDPL
constant Tile_X22Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000001010101000000000101010100000000000000000000000001010101000000000101010101010101000000000000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000111111111111111101000100010001000000000000000000";
--X23Y53, linear_LMDPL
constant Tile_X23Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000000000000000000000000000010101010000000010101010000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X24Y53, nonlinear_LMDPL
constant Tile_X24Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101101010100000000000000000000000001010101010101010010101010000000000000000000000000000000000000000101010101010101010101010010001000100010000000000101010100000000000000000101010101010101011011101110111010000000000000000";
--X25Y53, linear_LMDPL
constant Tile_X25Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000111111110000000010101010010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X26Y53, linear_LMDPL
constant Tile_X26Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010010101010101010100000000000000001111111111111111000000000000000011101110111011100000000000000000";
--X27Y53, nonlinear_LMDPL
constant Tile_X27Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111110101010010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X28Y53, linear_LMDPL
constant Tile_X28Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000101010101010101000000000000000000000000000000001010101010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001000100010001000";
--X29Y53, linear_LMDPL
constant Tile_X29Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010101010101000000001010101000000000000000001010101010101010010101010101010100000000000000000000000000000000000000000000000010111011101110110000000000000000";
--X30Y53, nonlinear_LMDPL
constant Tile_X30Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X31Y53, linear_LMDPL
constant Tile_X31Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000001010101010101010010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X32Y53, linear_LMDPL
constant Tile_X32Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010111111110000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000111011101110111000000000000000001000100010001000000000000000000";
--X33Y53, nonlinear_LMDPL
constant Tile_X33Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000011111111000000001010101000000000101010100000000000000000000100010001000100000000010101010010001000100010000000000000000000000000000000000100010001000100";
--X34Y53, linear_LMDPL
constant Tile_X34Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X35Y53, linear_LMDPL
constant Tile_X35Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000001010101010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X36Y53, nonlinear_LMDPL
constant Tile_X36Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010010101010000000010101010000000001010101000000000101010101010101001010101010001000100010000000000101010100000000000000000010001000100010001000100010001000000000000000000";
--X37Y53, linear_LMDPL
constant Tile_X37Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101111111110000000010101010010101010101010100000000000000001110111011101110000000000000000010111011101110110000000000000000";
--X38Y53, linear_LMDPL
constant Tile_X38Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X39Y53, nonlinear_LMDPL
constant Tile_X39Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000001010101001010101101010100000000011111111010101010101010100000000101010100010001000100010000000000000000010101010101010100000000000000000";
--X40Y53, linear_LMDPL
constant Tile_X40Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000101010101010101";
--X41Y53, linear_LMDPL
constant Tile_X41Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000101010100000000001010101010101010101010100000000101010101000100010001000000000000000000010101010101010100000000000000000";
--X42Y53, nonlinear_LMDPL
constant Tile_X42Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000101110111011101100000000000000000010001000100010";
--X43Y53, linear_LMDPL
constant Tile_X43Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000001010101101010100000000010101010000000001010101011111111010101010000000010101010000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101010111011101110110000000000000000";
--X44Y53, linear_LMDPL
constant Tile_X44Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010110101010010101010000000000000000101010100000000000000000111111110000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000011001100110011001100110011001100000000000000000";
--X45Y53, nonlinear_LMDPL
constant Tile_X45Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101010101010101010100101010100000000000000000000000000000000000000000000000011111111000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X46Y53, linear_LMDPL
constant Tile_X46Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000101010110101010000000000000000011111111000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X47Y53, linear_LMDPL
constant Tile_X47Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X48Y53, nonlinear_LMDPL
constant Tile_X48Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X49Y53, linear_LMDPL
constant Tile_X49Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000000000000000000011111111111111110000000000000000";
--X50Y53, linear_LMDPL
constant Tile_X50Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000010101010101010100000000010101010010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X51Y53, nonlinear_LMDPL
constant Tile_X51Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110101010110101010000000001010101000000000000000000000000010101010010101010101010100000000101010100000000000000000000000000000000010111011101110110000000000000000";
--X52Y53, linear_LMDPL
constant Tile_X52Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000001000100010001001100110011001100000000000000000";
--X53Y53, linear_LMDPL
constant Tile_X53Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000101010100000000000000001010101000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X54Y53, nonlinear_LMDPL
constant Tile_X54Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101110111011101110110000000000000000";
--X55Y53, linear_LMDPL
constant Tile_X55Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101011111111000000000000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000101010101010101001000100010001000000000000000000";
--X56Y53, linear_LMDPL
constant Tile_X56Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001111111111111111";
--X57Y53, nonlinear_LMDPL
constant Tile_X57Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X58Y53, linear_LMDPL
constant Tile_X58Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010101010101010100000000000000001110111011101110";
--X59Y53, linear_LMDPL
constant Tile_X59Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111101010101010101010101010111111111101010101100110011001100000000000000000000100010001000100000000000000000";
--X60Y53, nonlinear_LMDPL
constant Tile_X60Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000001010101010101010000000000000000000000000000000000101010110101010101010100000000010101010000000000000000000000000000000000000000010101010010001000100010000000000101010100000000000000000100010001000100000000000000000000000000000000000";
--X61Y53, linear_LMDPL
constant Tile_X61Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X62Y53, linear_LMDPL
constant Tile_X62Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000000110011001100110";
--X63Y53, nonlinear_LMDPL
constant Tile_X63Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000101010100000000010101010000100010001000100000000101010100010001000100010000000000000000000000000000000001010101010101010";
--X64Y53, linear_LMDPL
constant Tile_X64Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000001010101001010101101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100100110011001100110000000000000000";
--X65Y53, linear_LMDPL
constant Tile_X65Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000010101010000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X66Y53, nonlinear_LMDPL
constant Tile_X66Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000000000000000000010101010000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X67Y53, linear_LMDPL
constant Tile_X67Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X68Y53, linear_LMDPL
constant Tile_X68Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101010101010000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000010101010000000000000000000000000000000000000000101010100000000010101010000100010001000110101010000000001100110011001100000000000000000000000000000000001101110111011101";
--X69Y53, nonlinear_LMDPL
constant Tile_X69Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000101010101010101000000000000000001000100010001000000000000000000";
--X70Y53, linear_LMDPL
constant Tile_X70Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010101010101010100100010001000100000000000000000";
--X71Y53, linear_LMDPL
constant Tile_X71Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000000011001100110011";
--X72Y53, nonlinear_LMDPL
constant Tile_X72Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000101010100000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X73Y53, linear_LMDPL
constant Tile_X73Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000001111111100000000000000000000000010101010010101010000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001100110011001100";
--X74Y53, linear_LMDPL
constant Tile_X74Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X75Y53, nonlinear_LMDPL
constant Tile_X75Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000011001100110011000000000000000000011001100110011";
--X76Y53, linear_LMDPL
constant Tile_X76Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X77Y53, linear_LMDPL
constant Tile_X77Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X78Y53, ctrl_to_sec
constant Tile_X78Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y53, combined_WDDL
constant Tile_X79Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y53, combined_WDDL
constant Tile_X80Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y53, ctrl_IO
constant Tile_X81Y53_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y54, W_IO_custom
constant Tile_X0Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000";
--X1Y54, linear_LMDPL
constant Tile_X1Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000101010110101010000100010001000100000000111111111100110011001100000000000000000000000000000000000100010001000100";
--X2Y54, linear_LMDPL
constant Tile_X2Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000010101010101010100000000000000001001100110011001000000000000000000110011001100110000000000000000";
--X3Y54, nonlinear_LMDPL
constant Tile_X3Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X4Y54, linear_LMDPL
constant Tile_X4Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010111111111010101000000000010101010101010100000000000000000010001000100010000000000000000010011001100110010000000000000000";
--X5Y54, linear_LMDPL
constant Tile_X5Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000101010100000000000000000000000000000000000000000000000001010101001010101010001000100010000000000000000000000000000000000101010101010101010011001100110010000000000000000";
--X6Y54, nonlinear_LMDPL
constant Tile_X6Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000110011001100110";
--X7Y54, linear_LMDPL
constant Tile_X7Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X8Y54, linear_LMDPL
constant Tile_X8Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000010101011111111100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X9Y54, nonlinear_LMDPL
constant Tile_X9Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X10Y54, linear_LMDPL
constant Tile_X10Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000001010101010101010010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X11Y54, linear_LMDPL
constant Tile_X11Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X12Y54, nonlinear_LMDPL
constant Tile_X12Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000001010101000000000000000001010101010101010010001000100010000000000000000000000000000000000101110111011101100010001000100010000000000000000";
--X13Y54, linear_LMDPL
constant Tile_X13Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000001010101010101010111111110000000000000000010101010101010100000000000000001001100110011001000000000000000010001000100010000000000000000000";
--X14Y54, linear_LMDPL
constant Tile_X14Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000010101010000000000000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X15Y54, nonlinear_LMDPL
constant Tile_X15Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000011001100110011";
--X16Y54, linear_LMDPL
constant Tile_X16Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000000100010001000100000000000000000000000000000000000000000000000000";
--X17Y54, linear_LMDPL
constant Tile_X17Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001000100010001000";
--X18Y54, nonlinear_LMDPL
constant Tile_X18Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000101010101010101000000000000000000111011101110111";
--X19Y54, linear_LMDPL
constant Tile_X19Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000111111110000000000000000000100010001000100000000101010101011101110111011000000000000000000000000000000001100110011001100";
--X20Y54, linear_LMDPL
constant Tile_X20Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X21Y54, nonlinear_LMDPL
constant Tile_X21Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000010101010101010100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000110011001100110000000000000000001101110111011101";
--X22Y54, linear_LMDPL
constant Tile_X22Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000001010101101010100000000000000000000000001010101000000000101010100000000011111111101010100000000000000000000000001010101010101010010101010101010100000000000000000110011001100110000000000000000000110011001100110000000000000000";
--X23Y54, linear_LMDPL
constant Tile_X23Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101011111111000000000101010101010101000000000000000000000000101010100000000000000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X24Y54, nonlinear_LMDPL
constant Tile_X24Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000011111111000000001010101010101010010101010000000000000000000000001010101000000000101010101010101000000000010001000100010000000000000000000000000000000000101110111011101110101010101010100000000000000000";
--X25Y54, linear_LMDPL
constant Tile_X25Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010101111111110101010010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X26Y54, linear_LMDPL
constant Tile_X26Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001111111100000000010101010101010100000000010101010110011001100110000000000000000011001100110011000000000000000000";
--X27Y54, nonlinear_LMDPL
constant Tile_X27Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001000100010001000";
--X28Y54, linear_LMDPL
constant Tile_X28Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001010101011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X29Y54, linear_LMDPL
constant Tile_X29Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000010101010000000001010101101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010010101010101010110101010101010101000100010001000000000000000000000000000000000000000000000000000";
--X30Y54, nonlinear_LMDPL
constant Tile_X30Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001101110111011101";
--X31Y54, linear_LMDPL
constant Tile_X31Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001011101110111011";
--X32Y54, linear_LMDPL
constant Tile_X32Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000101010110101010000000001111111100000000000000000000000000000000000100010001000110101010000000000010001000100010000000000000000000000000000000000000000000000000";
--X33Y54, nonlinear_LMDPL
constant Tile_X33Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111110101010000000000000000000000000000000001010101010101010101010100000000000000000000000001010101000000000101010100000000000000000010101010101010100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X34Y54, linear_LMDPL
constant Tile_X34Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000100010001000100000000000000000000110011001100110000000000000000";
--X35Y54, linear_LMDPL
constant Tile_X35Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010100000000010101010000100010001000111111111000000000101010101010101000000000000000000000000000000000000000000000000";
--X36Y54, nonlinear_LMDPL
constant Tile_X36Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000101010110101010000000001010101000000000000000000000000011111111010101010101010100000000101010101011101110111011000000000000000010101010101010100000000000000000";
--X37Y54, linear_LMDPL
constant Tile_X37Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010101010110101010000000001100110011001100000000000000000010111011101110110000000000000000";
--X38Y54, linear_LMDPL
constant Tile_X38Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000010101010101010100000000101010100000000000000000000000000000000011001100110011000000000000000000";
--X39Y54, nonlinear_LMDPL
constant Tile_X39Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000000000000010101010000100010001000100000000101010101100110011001100000000000000000000000000000000001101110111011101";
--X40Y54, linear_LMDPL
constant Tile_X40Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000011111111010101010101010100000000111111111110111011101110000000000000000001000100010001000000000000000000";
--X41Y54, linear_LMDPL
constant Tile_X41Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010111111111101010101010101010101010000000000000000001000100010001000000000000000000";
--X42Y54, nonlinear_LMDPL
constant Tile_X42Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010101010000000010101010010101011010101010101010000000001010101010101010000000000000000010101010000100010001000100000000101010100101010101010101000000000000000000000000000000000110011001100110";
--X43Y54, linear_LMDPL
constant Tile_X43Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000101010100000000000000000000000010101010000000001010101000000000101010100000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X44Y54, linear_LMDPL
constant Tile_X44Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000010101010000000000000000000000000000000000000000000000000010101010101010110101010000000000000000010101010101010100000000010101010000000000000000000000000000000000000000000000000101110111011101100000000000000001100110011001100";
--X45Y54, nonlinear_LMDPL
constant Tile_X45Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010111111110101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000110011001100110";
--X46Y54, linear_LMDPL
constant Tile_X46Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000000000001111111100000000010101011010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X47Y54, linear_LMDPL
constant Tile_X47Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010110101010000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000100010001000100010111011101110110000000000000000";
--X48Y54, nonlinear_LMDPL
constant Tile_X48Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X49Y54, linear_LMDPL
constant Tile_X49Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010101010100101010111111111010101010101010100000000101010101100110011001100000000000000000011101110111011100000000000000000";
--X50Y54, linear_LMDPL
constant Tile_X50Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111110101010000000001010101010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000010101010101010110101010000000001000100010001000000000000000000000100010001000100000000000000000";
--X51Y54, nonlinear_LMDPL
constant Tile_X51Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101001010101101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000000000000111111110101010110101010000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000000000100010001000100000000000000000000011001100110011";
--X52Y54, linear_LMDPL
constant Tile_X52Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000010001000100010000000000000000000000000000000000001100110011001110111011101110110000000000000000";
--X53Y54, linear_LMDPL
constant Tile_X53Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000111111110000000000000000010101010101010110111011101110110000000000000000";
--X54Y54, nonlinear_LMDPL
constant Tile_X54Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X55Y54, linear_LMDPL
constant Tile_X55Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010101010101000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001000100010001000";
--X56Y54, linear_LMDPL
constant Tile_X56Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001010101010101010";
--X57Y54, nonlinear_LMDPL
constant Tile_X57Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000110011001100110";
--X58Y54, linear_LMDPL
constant Tile_X58Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000001010101001010101000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X59Y54, linear_LMDPL
constant Tile_X59Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101001010101010001000100010010101010111111110000000000000000001000100010001010101010101010100000000000000000";
--X60Y54, nonlinear_LMDPL
constant Tile_X60Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000010101010101010100000000010101010000000001010101000000000000000001010101010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X61Y54, linear_LMDPL
constant Tile_X61Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000001111111100000000111111110000000000000000101010100000000010101010000000000000000011111111000000000000000000000000000000000000000010101010010101010101010110101010000000001100110011001100000000000000000011111111111111110000000000000000";
--X62Y54, linear_LMDPL
constant Tile_X62Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000001010101000000000000000000000000011111111000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000010001000100010001000100010001000000000000000000";
--X63Y54, nonlinear_LMDPL
constant Tile_X63Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000010101010010101010000000010101010000000001010101000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X64Y54, linear_LMDPL
constant Tile_X64Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000010001000100010000000000000000000000000000000000011001100110011";
--X65Y54, linear_LMDPL
constant Tile_X65Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110111011101110110001000100010000000000000000000";
--X66Y54, nonlinear_LMDPL
constant Tile_X66Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000010001000100010000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X67Y54, linear_LMDPL
constant Tile_X67Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000001000100010001000";
--X68Y54, linear_LMDPL
constant Tile_X68Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000001111111111111111";
--X69Y54, nonlinear_LMDPL
constant Tile_X69Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y54, linear_LMDPL
constant Tile_X70Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001111111100000000000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000000010001000100010";
--X71Y54, linear_LMDPL
constant Tile_X71Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000001010101011111111000000000000000000000000010101010000000000000000010101010101010100000000000000001101110111011101000000000000000010101010101010100000000000000000";
--X72Y54, nonlinear_LMDPL
constant Tile_X72Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000010101010000000000000000010101010101010100000000000000000001000100010001000000000000000001000100010001000000000000000000";
--X73Y54, linear_LMDPL
constant Tile_X73Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000000000000001000100010001000000000000000000000000000000000100010001000100";
--X74Y54, linear_LMDPL
constant Tile_X74Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111101010100000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001010101010101010";
--X75Y54, nonlinear_LMDPL
constant Tile_X75Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X76Y54, linear_LMDPL
constant Tile_X76Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010011001100110010000000000000000";
--X77Y54, linear_LMDPL
constant Tile_X77Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000001000100010001";
--X78Y54, ctrl_to_sec
constant Tile_X78Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y54, combined_WDDL
constant Tile_X79Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y54, combined_WDDL
constant Tile_X80Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y54, ctrl_IO
constant Tile_X81Y54_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y55, W_IO_custom
constant Tile_X0Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000";
--X1Y55, linear_LMDPL
constant Tile_X1Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000010101010101010100000000000000001111111111111111000000000000000010101010101010100000000000000000";
--X2Y55, linear_LMDPL
constant Tile_X2Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000010101010010101010000000000000000010001000100010000000000101010100000000000000000001000100010001010111011101110110000000000000000";
--X3Y55, nonlinear_LMDPL
constant Tile_X3Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000010001000100010000000000000000000010001000100010000000000000000";
--X4Y55, linear_LMDPL
constant Tile_X4Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000010101010000000001111111100000000101010101010101000000000010001000100010000000000000000000000000000000000001100110011001110111011101110110000000000000000";
--X5Y55, linear_LMDPL
constant Tile_X5Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X6Y55, nonlinear_LMDPL
constant Tile_X6Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000000000000000000";
--X7Y55, linear_LMDPL
constant Tile_X7Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X8Y55, linear_LMDPL
constant Tile_X8Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X9Y55, nonlinear_LMDPL
constant Tile_X9Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110011001100110000000000000000000011001100110011";
--X10Y55, linear_LMDPL
constant Tile_X10Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001001100110011001";
--X11Y55, linear_LMDPL
constant Tile_X11Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010010101010101010100000000000000000010001000100010000000000000000010101010101010100000000000000000";
--X12Y55, nonlinear_LMDPL
constant Tile_X12Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000010101010000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001100110011001100";
--X13Y55, linear_LMDPL
constant Tile_X13Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000101010100000000000000000000000000101010110101010000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000000100010001000111001100110011000000000000000000";
--X14Y55, linear_LMDPL
constant Tile_X14Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000001010101000000000000000000000000000000000000000000000000010101010101010101010101101010101000100010001000000000000000000010101010101010100000000000000000";
--X15Y55, nonlinear_LMDPL
constant Tile_X15Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001010101000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000100110011001100100000000000000000011001100110011";
--X16Y55, linear_LMDPL
constant Tile_X16Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000110101010000000001011101110111011000000000000000000000000000000000011001100110011";
--X17Y55, linear_LMDPL
constant Tile_X17Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010000000000000000000000000000001010101011111111010101010000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X18Y55, nonlinear_LMDPL
constant Tile_X18Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110101010101010101000000001010101010101010010101010000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X19Y55, linear_LMDPL
constant Tile_X19Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010110101010000000000000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000011101110111011111001100110011000000000000000000";
--X20Y55, linear_LMDPL
constant Tile_X20Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100011001100110011000000000000000000";
--X21Y55, nonlinear_LMDPL
constant Tile_X21Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100101010101010101000000001010101000000000000000000101010100000000010001000100010000000000101010100000000000000000001100110011001110011001100110010000000000000000";
--X22Y55, linear_LMDPL
constant Tile_X22Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000001010101010101010101010100101010100000000111111110000000000000000000000000000000010101010010101010101010110101010000000001000100010001000000000000000000001000100010001000000000000000000";
--X23Y55, linear_LMDPL
constant Tile_X23Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101011010101000000000000000000000000001010101000000000000000001010101010101010000000000000000111111110000000000000000000000001010101000000000000000000000000000000000101010100101010100000000000100010001000100000000000000000100010001000100000000000000000000000000000000001101110111011101";
--X24Y55, nonlinear_LMDPL
constant Tile_X24Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101010101000000000010101010101010100000000101010101010101010101010000000000000000000100010001000100000000000000000";
--X25Y55, linear_LMDPL
constant Tile_X25Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000101010100101010110101010000100010001000100000000000000001011101110111011000000000000000000000000000000000010001000100010";
--X26Y55, linear_LMDPL
constant Tile_X26Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100110011001100110000000000000000";
--X27Y55, nonlinear_LMDPL
constant Tile_X27Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000001010101010101010010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X28Y55, linear_LMDPL
constant Tile_X28Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000010101010010101010000000000000000101010100000000000000000000000000101010100000000000000000000000000000000000000001010101000000000010101010101010100000000111111111010101010101010000000000000000011111111111111110000000000000000";
--X29Y55, linear_LMDPL
constant Tile_X29Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000001010101010101010010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X30Y55, nonlinear_LMDPL
constant Tile_X30Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000011111111000000000000000000000000000000000000000000000000011001100110011000000000000000001011101110111011";
--X31Y55, linear_LMDPL
constant Tile_X31Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001100110011001100";
--X32Y55, linear_LMDPL
constant Tile_X32Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000101010110101010000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000010101010101010100000000000000001111111111111111";
--X33Y55, nonlinear_LMDPL
constant Tile_X33Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101010101010101010100000000000000000000000001010101000000000000000000000000001010101000100010001000100000000101010101100110011001100000000000000000000000000000000000100010001000100";
--X34Y55, linear_LMDPL
constant Tile_X34Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000001010101011111111000000000000000000000000000000000000000000000000010101010101010100000000010101010000000000000000000000000000000001100110011001100000000000000000";
--X35Y55, linear_LMDPL
constant Tile_X35Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000010101010000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X36Y55, nonlinear_LMDPL
constant Tile_X36Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000010101010000000001010101000000000000000001010101000000000000000000000000010101010010001000100010000000000101010100000000000000000001000100010001010001000100010000000000000000000";
--X37Y55, linear_LMDPL
constant Tile_X37Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000010101010000000000000000010101010010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X38Y55, linear_LMDPL
constant Tile_X38Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000000001010101000000000000000001111111100000000000100010001000100000000000000001011101110111011000000000000000000000000000000000011001100110011";
--X39Y55, nonlinear_LMDPL
constant Tile_X39Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000011111111010101010101010100000000101010101000100010001000000000000000000000000000000000000000000000000000";
--X40Y55, linear_LMDPL
constant Tile_X40Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000010101010000000000000000011111111000000000000000000000000001000100010001000000000000000000000000000000000";
--X41Y55, linear_LMDPL
constant Tile_X41Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000010101010010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X42Y55, nonlinear_LMDPL
constant Tile_X42Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101010101010000000000000000000000000101010100000000010101010000100010001000100000000101010100000000000000000000000000000000000000000000000001101110111011101";
--X43Y55, linear_LMDPL
constant Tile_X43Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010110101010000000000000000010101010000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000101010101010101000000000000000000100010001000100";
--X44Y55, linear_LMDPL
constant Tile_X44Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101010101010000000000101010100000000000000000000000000000000101010101111111100000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X45Y55, nonlinear_LMDPL
constant Tile_X45Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X46Y55, linear_LMDPL
constant Tile_X46Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000101010100101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000010001000100010";
--X47Y55, linear_LMDPL
constant Tile_X47Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X48Y55, nonlinear_LMDPL
constant Tile_X48Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000111111110000000000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X49Y55, linear_LMDPL
constant Tile_X49Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000111111111010101010101010010101010101010100000000000000000010001000100010000000000000000011001100110011000000000000000000";
--X50Y55, linear_LMDPL
constant Tile_X50Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000010001000100010000000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X51Y55, nonlinear_LMDPL
constant Tile_X51Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001111111100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010101010101010101010000000001010101001010101101010101010101010101010010101010101010100000000101010100011001100110011000000000000000011001100110011000000000000000000";
--X52Y55, linear_LMDPL
constant Tile_X52Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X53Y55, linear_LMDPL
constant Tile_X53Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000011111111000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001100110011001100";
--X54Y55, nonlinear_LMDPL
constant Tile_X54Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X55Y55, linear_LMDPL
constant Tile_X55Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000010101010101010100000000000000000000000001111111100000000101010100000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X56Y55, linear_LMDPL
constant Tile_X56Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001000100010001000";
--X57Y55, nonlinear_LMDPL
constant Tile_X57Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000110011001100110000000000000000000100010001000100";
--X58Y55, linear_LMDPL
constant Tile_X58Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000000000001010101010101010000000000000000000000000010101010000000000000000001000100010001000000000000000000001000100010001";
--X59Y55, linear_LMDPL
constant Tile_X59Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X60Y55, nonlinear_LMDPL
constant Tile_X60Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000010101010010101010000000010101010000000000000000000000000000000000000000001010101000100010001000100000000101010100000000000000000000000000000000000000000000000000001000100010001";
--X61Y55, linear_LMDPL
constant Tile_X61Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111111111111100000000000000000010001000100010";
--X62Y55, linear_LMDPL
constant Tile_X62Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000111111110000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001010101010101010";
--X63Y55, nonlinear_LMDPL
constant Tile_X63Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010010101010000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000101010100100010001000100000000000000000000000000000000001100110011001100";
--X64Y55, linear_LMDPL
constant Tile_X64Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000001010101000000000000000010101010101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X65Y55, linear_LMDPL
constant Tile_X65Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000101010100000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X66Y55, nonlinear_LMDPL
constant Tile_X66Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000001010101000000000101010100000000000000000010001000100010000000000000000000000000000000000000100010001000100110011001100110000000000000000";
--X67Y55, linear_LMDPL
constant Tile_X67Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000100010001000100";
--X68Y55, linear_LMDPL
constant Tile_X68Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010110101010000000001100110011001100000000000000000010101010101010100000000000000000";
--X69Y55, nonlinear_LMDPL
constant Tile_X69Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010100000000000000000000000000000000000000000111111110000000010101010000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X70Y55, linear_LMDPL
constant Tile_X70Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X71Y55, linear_LMDPL
constant Tile_X71Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X72Y55, nonlinear_LMDPL
constant Tile_X72Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000001010101010101010000000001010101000000000101010101111111100000000010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X73Y55, linear_LMDPL
constant Tile_X73Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000001000100010001";
--X74Y55, linear_LMDPL
constant Tile_X74Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000011001100110011";
--X75Y55, nonlinear_LMDPL
constant Tile_X75Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X76Y55, linear_LMDPL
constant Tile_X76Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000011001100110011";
--X77Y55, linear_LMDPL
constant Tile_X77Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001001100110011001000000000000000010001000100010000000000000000000";
--X78Y55, ctrl_to_sec
constant Tile_X78Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y55, combined_WDDL
constant Tile_X79Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y55, combined_WDDL
constant Tile_X80Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y55, ctrl_IO
constant Tile_X81Y55_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y56, W_IO_custom
constant Tile_X0Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y56, linear_LMDPL
constant Tile_X1Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000111111111010101000000000010001000100010000000000000000000000000000000000001100110011001111101110111011100000000000000000";
--X2Y56, linear_LMDPL
constant Tile_X2Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010101010101010100000000000000001001100110011001000000000000000011001100110011000000000000000000";
--X3Y56, nonlinear_LMDPL
constant Tile_X3Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010101010100000000000000000100010001000100000000000000000000110011001100110000000000000000";
--X4Y56, linear_LMDPL
constant Tile_X4Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000010101010101010101010101000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X5Y56, linear_LMDPL
constant Tile_X5Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000001101110111011101";
--X6Y56, nonlinear_LMDPL
constant Tile_X6Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X7Y56, linear_LMDPL
constant Tile_X7Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001000100010001000000000000000000011111111111111110000000000000000";
--X8Y56, linear_LMDPL
constant Tile_X8Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X9Y56, nonlinear_LMDPL
constant Tile_X9Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X10Y56, linear_LMDPL
constant Tile_X10Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X11Y56, linear_LMDPL
constant Tile_X11Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010010101010101010100000000000000000000000000000000000000000000000011001100110011000000000000000000";
--X12Y56, nonlinear_LMDPL
constant Tile_X12Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010101010100000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010100001000100010001000000000000000010001000100010000000000000000000";
--X13Y56, linear_LMDPL
constant Tile_X13Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000001000100010001000";
--X14Y56, linear_LMDPL
constant Tile_X14Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X15Y56, nonlinear_LMDPL
constant Tile_X15Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000101010100000000101010100000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000110111011101110111001100110011000000000000000000";
--X16Y56, linear_LMDPL
constant Tile_X16Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001111111111111111000000000000000000000000000000000100010001000100";
--X17Y56, linear_LMDPL
constant Tile_X17Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X18Y56, nonlinear_LMDPL
constant Tile_X18Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000001010101010101010000000001010101000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X19Y56, linear_LMDPL
constant Tile_X19Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000101010101011101110111011000000000000000011001100110011000000000000000000";
--X20Y56, linear_LMDPL
constant Tile_X20Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X21Y56, nonlinear_LMDPL
constant Tile_X21Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111111010101010101010101010100000000010101010000000001010101000000000000000001010101001010101000100010001000100000000101010100001000100010001000000000000000000000000000000001000100010001000";
--X22Y56, linear_LMDPL
constant Tile_X22Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000001010101010101010111111110000000000000000111111110000000000000000000000000000000010101010010101010101010100000000000000000101010101010101000000000000000001000100010001000000000000000000";
--X23Y56, linear_LMDPL
constant Tile_X23Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100101010100000000000000000000000001010101000000000000000010101010000000000000000000000000000000001010101000000000000000000101010101010101000000000000000000000000101010101010101000000000010101010101010100000000000000000011001100110011000000000000000001110111011101110000000000000000";
--X24Y56, nonlinear_LMDPL
constant Tile_X24Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010101010101000000000010001000100010000000000010101010000000000000000100010001000100001000100010001000000000000000000";
--X25Y56, linear_LMDPL
constant Tile_X25Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000101010101010101011111111000000000000000000000000101010101111111100000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X26Y56, linear_LMDPL
constant Tile_X26Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000001111111100000000000000000000000010101010000000000000000010101010000000000000000000000000000100010001000100000000000000000101010101010101000000000000000000000000000000001010101010101010";
--X27Y56, nonlinear_LMDPL
constant Tile_X27Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001100110011001110001000100010000000000000000000";
--X28Y56, linear_LMDPL
constant Tile_X28Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001010101011111111000100010001000100000000000000001100110011001100000000000000000000000000000000000011001100110011";
--X29Y56, linear_LMDPL
constant Tile_X29Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000010101010000000000101010111111111000000000000000000000000000000001010101010101010000100010001000100000000101010100000000000000000000000000000000000000000000000001110111011101110";
--X30Y56, nonlinear_LMDPL
constant Tile_X30Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X31Y56, linear_LMDPL
constant Tile_X31Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111110101010000000000000000011111111000000000000000000000000000000001010101010101010010001000100010000000000000000000000000000000000111011101110111000000000000000000000000000000000";
--X32Y56, linear_LMDPL
constant Tile_X32Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000010101010010101010101010100000000010101010100010001000100000000000000000000110011001100110000000000000000";
--X33Y56, nonlinear_LMDPL
constant Tile_X33Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000010101010101010100101010100000000000000001010101000000000101010100000000010101010010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X34Y56, linear_LMDPL
constant Tile_X34Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X35Y56, linear_LMDPL
constant Tile_X35Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000000000101010100000000000000000000000011111111101010100000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X36Y56, nonlinear_LMDPL
constant Tile_X36Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000010101010000000001010101011111111000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000001100110011001100000000000000001100110011001100";
--X37Y56, linear_LMDPL
constant Tile_X37Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X38Y56, linear_LMDPL
constant Tile_X38Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000101010100000000000000000000000011111111000000001111111100000000000100010001000100000000010101011011101110111011000000000000000000000000000000000100010001000100";
--X39Y56, nonlinear_LMDPL
constant Tile_X39Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000001010101000000000111111110000000000000000010101010101010100000000101010100100010001000100000000000000000000100010001000100000000000000000";
--X40Y56, linear_LMDPL
constant Tile_X40Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101010101010101010100000000000000001100110011001100000000000000000011101110111011100000000000000000";
--X41Y56, linear_LMDPL
constant Tile_X41Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010000100010001000100000000101010101000100010001000000000000000000000000000000000000010001000100010";
--X42Y56, nonlinear_LMDPL
constant Tile_X42Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000010101010000000001010101010101010111111110000000010101010010101010101010100000000000000001101110111011101000000000000000011001100110011000000000000000000";
--X43Y56, linear_LMDPL
constant Tile_X43Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000001111111100000000101010100000000010101010010101010101010100000000000000000100010001000100000000000000000010001000100010000000000000000000";
--X44Y56, linear_LMDPL
constant Tile_X44Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000000000000001010101000000000000000000000000010101011010101010101010000000000000000000000000000000000000000010101010111111110000000000000000010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X45Y56, nonlinear_LMDPL
constant Tile_X45Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000001010101010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X46Y56, linear_LMDPL
constant Tile_X46Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001011101110111011";
--X47Y56, linear_LMDPL
constant Tile_X47Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001010101010101010";
--X48Y56, nonlinear_LMDPL
constant Tile_X48Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000011111111010101010101010100000000101010100100010001000100000000000000000000100010001000100000000000000000";
--X49Y56, linear_LMDPL
constant Tile_X49Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000010101010101010100000000000000001110111011101110000000000000000011001100110011000000000000000000";
--X50Y56, linear_LMDPL
constant Tile_X50Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000101010101010101011111111000100010001000100000000000000000010001000100010000000000000000000000000000000000000000000000000";
--X51Y56, nonlinear_LMDPL
constant Tile_X51Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000111111111010101010101010000000001010101000000000000000001010101000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000011001100110011";
--X52Y56, linear_LMDPL
constant Tile_X52Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X53Y56, linear_LMDPL
constant Tile_X53Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100000000000000000000000000000000000110011001100110000000000000000";
--X54Y56, nonlinear_LMDPL
constant Tile_X54Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X55Y56, linear_LMDPL
constant Tile_X55Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X56Y56, linear_LMDPL
constant Tile_X56Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001000100010001000000000000000000";
--X57Y56, nonlinear_LMDPL
constant Tile_X57Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X58Y56, linear_LMDPL
constant Tile_X58Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X59Y56, linear_LMDPL
constant Tile_X59Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010010101010101010110101010000000001010101010101010000000000000000011101110111011100000000000000000";
--X60Y56, nonlinear_LMDPL
constant Tile_X60Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000000000000000000011111111000100010001000100000000000000001010101010101010000000000000000000000000000000000001000100010001";
--X61Y56, linear_LMDPL
constant Tile_X61Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000101010100000000010101010010001000100010000000000000000000000000000000000101010101010101001100110011001100000000000000000";
--X62Y56, linear_LMDPL
constant Tile_X62Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000011111111010101010101010100000000000000001101110111011101000000000000000010111011101110110000000000000000";
--X63Y56, nonlinear_LMDPL
constant Tile_X63Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000010101010000000001010101000000000000000000000000010101010000100010001000100000000000000000011001100110011000000000000000000000000000000000000000000000000";
--X64Y56, linear_LMDPL
constant Tile_X64Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000001111111101010101101010100000000000000000000000000000000000000000000000000000000001010101010001000100010000000000000000000000000000000000100010001000100000100010001000100000000000000000";
--X65Y56, linear_LMDPL
constant Tile_X65Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X66Y56, nonlinear_LMDPL
constant Tile_X66Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000001010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000000100010001000100";
--X67Y56, linear_LMDPL
constant Tile_X67Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000011001100110011000000000000000000001000100010001";
--X68Y56, linear_LMDPL
constant Tile_X68Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001111111111111111000000000000000010101010101010100000000000000000";
--X69Y56, nonlinear_LMDPL
constant Tile_X69Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000010101010000000000000000010101010000100010001000100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X70Y56, linear_LMDPL
constant Tile_X70Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X71Y56, linear_LMDPL
constant Tile_X71Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X72Y56, nonlinear_LMDPL
constant Tile_X72Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010101010101000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000100010001000100";
--X73Y56, linear_LMDPL
constant Tile_X73Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X74Y56, linear_LMDPL
constant Tile_X74Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000101010101010101";
--X75Y56, nonlinear_LMDPL
constant Tile_X75Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000000000000101010100000000000000000000000000000000010101010000000000000000010101010101010100000000000000000100010001000100000000000000000000010001000100010000000000000000";
--X76Y56, linear_LMDPL
constant Tile_X76Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000100010001000100000000000000001011101110111011000000000000000000000000000000000111011101110111";
--X77Y56, linear_LMDPL
constant Tile_X77Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000111111111010101010101010000000000000000000000000000000000000000000000000";
--X78Y56, ctrl_to_sec
constant Tile_X78Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y56, combined_WDDL
constant Tile_X79Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y56, combined_WDDL
constant Tile_X80Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y56, ctrl_IO
constant Tile_X81Y56_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y57, W_IO_custom
constant Tile_X0Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y57, linear_LMDPL
constant Tile_X1Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001111111100000000010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X2Y57, linear_LMDPL
constant Tile_X2Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111110101010000000000000000000000000101010100000000000000000010101010101010100000000000000001101110111011101000000000000000011101110111011100000000000000000";
--X3Y57, nonlinear_LMDPL
constant Tile_X3Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000010101010010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X4Y57, linear_LMDPL
constant Tile_X4Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010101010100000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000100010001000100000000000000001100110011001100000000000000000000000000000000000110011001100110";
--X5Y57, linear_LMDPL
constant Tile_X5Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000001100110011001100";
--X6Y57, nonlinear_LMDPL
constant Tile_X6Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000010101010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001000100010001000";
--X7Y57, linear_LMDPL
constant Tile_X7Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000000110011001100110000000000000000";
--X8Y57, linear_LMDPL
constant Tile_X8Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001001100110011001000000000000000010111011101110110000000000000000";
--X9Y57, nonlinear_LMDPL
constant Tile_X9Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X10Y57, linear_LMDPL
constant Tile_X10Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000001000100010001000000000000000000";
--X11Y57, linear_LMDPL
constant Tile_X11Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010101011111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X12Y57, nonlinear_LMDPL
constant Tile_X12Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001001100110011001";
--X13Y57, linear_LMDPL
constant Tile_X13Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000101010101010101001000100010001000000000000000000";
--X14Y57, linear_LMDPL
constant Tile_X14Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000001010101001010101000000000000000001010101000000000000000000000000010001000100010000000000000000000000000000000000111111111111111101010101010101010000000000000000";
--X15Y57, nonlinear_LMDPL
constant Tile_X15Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000101010100000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000010001000100010";
--X16Y57, linear_LMDPL
constant Tile_X16Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000010001000100010000000000000000000000000000000000111111111111111110101010101010100000000000000000";
--X17Y57, linear_LMDPL
constant Tile_X17Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000001100110011001101000100010001000000000000000000";
--X18Y57, nonlinear_LMDPL
constant Tile_X18Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000001010101010101010000000000000000011111111000100010001000100000000000000001001100110011001000000000000000000000000000000001000100010001000";
--X19Y57, linear_LMDPL
constant Tile_X19Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000110011001100110";
--X20Y57, linear_LMDPL
constant Tile_X20Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000000011001100110011000000000000000001000100010001000000000000000000";
--X21Y57, nonlinear_LMDPL
constant Tile_X21Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000010101010000000000000000000000000000000010101010111111110000000010101010000000001010101000000000000000000101010101010101010001000100010000000000101010100000000000000000000000000000000000010001000100010000000000000000";
--X22Y57, linear_LMDPL
constant Tile_X22Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000101010110101010000000000000000000000000101010100000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X23Y57, linear_LMDPL
constant Tile_X23Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000001010101000000000101010110101010010101010000000000000000101010100000000000000000000000001010101011111111000000000000000000000000101010100000000000000000010101010101010100000000000000000010001000100010000000000000000010111011101110110000000000000000";
--X24Y57, nonlinear_LMDPL
constant Tile_X24Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000010101010101010100000000101010100100010001000100000000000000000000110011001100110000000000000000";
--X25Y57, linear_LMDPL
constant Tile_X25Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010101010100000000001010101000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X26Y57, linear_LMDPL
constant Tile_X26Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000000100010001000100000000000000001000100010001000000000000000000000000000000000001101110111011101";
--X27Y57, nonlinear_LMDPL
constant Tile_X27Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000011111111000000000000000000000000000000000000000001010101010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X28Y57, linear_LMDPL
constant Tile_X28Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000101010100000000000000000000000001111111110101010010101010000000000000000101010100000000000000000111111111010101011111111000000000000000000000000000000001010101010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000100010001000100";
--X29Y57, linear_LMDPL
constant Tile_X29Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000101010100000000000000001010101000000000010101011111111110101010010101010101010110101010000000001011101110111011000000000000000010001000100010000000000000000000";
--X30Y57, nonlinear_LMDPL
constant Tile_X30Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000110011001100110";
--X31Y57, linear_LMDPL
constant Tile_X31Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X32Y57, linear_LMDPL
constant Tile_X32Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000010101011010101001010101101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000100010001000110101010000000000010001000100010000000000000000000000000000000001010101010101010";
--X33Y57, nonlinear_LMDPL
constant Tile_X33Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000101010110101010101010101010101010101010000000001010101000000000101010100000000000000000000100010001000100000000101010101010101010101010000000000000000000000000000000001100110011001100";
--X34Y57, linear_LMDPL
constant Tile_X34Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000011101110111011100000000000000000";
--X35Y57, linear_LMDPL
constant Tile_X35Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010101010100000000000000001111111111111111000000000000000011001100110011000000000000000000";
--X36Y57, nonlinear_LMDPL
constant Tile_X36Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101010101010000000001010101000000000000000001010101011111111010001000100010000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X37Y57, linear_LMDPL
constant Tile_X37Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001111111100000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000100010001000110101010000000000100010001000100000000000000000000000000000000000010001000100010";
--X38Y57, linear_LMDPL
constant Tile_X38Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011";
--X39Y57, nonlinear_LMDPL
constant Tile_X39Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X40Y57, linear_LMDPL
constant Tile_X40Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000010001000100010010101010101010100000000000000000";
--X41Y57, linear_LMDPL
constant Tile_X41Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000001010101010101010101010100000000101010101111111111111111000000000000000011101110111011100000000000000000";
--X42Y57, nonlinear_LMDPL
constant Tile_X42Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101111111110000000010101010000000000000000000000000000000000000000010101010000100010001000100000000101010100011001100110011000000000000000000000000000000000000000000000000";
--X43Y57, linear_LMDPL
constant Tile_X43Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000001010101000000001010101000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001100110011001100000000000000000000000000000000000010001000100010";
--X44Y57, linear_LMDPL
constant Tile_X44Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000101010100101010110101010000000000101010100000000000000000000000000000000000000000000000011111111000100010001000100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X45Y57, nonlinear_LMDPL
constant Tile_X45Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X46Y57, linear_LMDPL
constant Tile_X46Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X47Y57, linear_LMDPL
constant Tile_X47Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000111111110000000001010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100000000000000000000000000000000001100110011001100";
--X48Y57, nonlinear_LMDPL
constant Tile_X48Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000001100110011001100000000000000001100110011001100";
--X49Y57, linear_LMDPL
constant Tile_X49Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X50Y57, linear_LMDPL
constant Tile_X50Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101011111111010101010101010100000000000000001011101110111011000000000000000011111111111111110000000000000000";
--X51Y57, nonlinear_LMDPL
constant Tile_X51Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000001010101000000000010001000100010000000000101010100000000000000000001000100010001011011101110111010000000000000000";
--X52Y57, linear_LMDPL
constant Tile_X52Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111000100010001000100000000000000001100110011001100000000000000000000000000000000000100010001000100";
--X53Y57, linear_LMDPL
constant Tile_X53Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000000000000000000011111111111111110000000000000000";
--X54Y57, nonlinear_LMDPL
constant Tile_X54Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000010101010000000000000000000000000000000000000000000000000000100010001000100000000000000000010001000100010000000000000000000000000000000000100010001000100";
--X55Y57, linear_LMDPL
constant Tile_X55Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000111011101110111000000000000000000000000000000001011101110111011";
--X56Y57, linear_LMDPL
constant Tile_X56Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000";
--X57Y57, nonlinear_LMDPL
constant Tile_X57Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000001010101010101010";
--X58Y57, linear_LMDPL
constant Tile_X58Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001011101110111011";
--X59Y57, linear_LMDPL
constant Tile_X59Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111111111110000000000000000010101010101010100000000000000001010101010101010000000000000000011111111111111110000000000000000";
--X60Y57, nonlinear_LMDPL
constant Tile_X60Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000100010001000100000000101010100011001100110011000000000000000000000000000000001001100110011001";
--X61Y57, linear_LMDPL
constant Tile_X61Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000101010100000000000000000010101010101010110101010000000001111111111111111000000000000000010101010101010100000000000000000";
--X62Y57, linear_LMDPL
constant Tile_X62Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001";
--X63Y57, nonlinear_LMDPL
constant Tile_X63Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000010001000100010000000000101010100000000000000000000100010001000110101010101010100000000000000000";
--X64Y57, linear_LMDPL
constant Tile_X64Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000000100010001000100000000000000000";
--X65Y57, linear_LMDPL
constant Tile_X65Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111110101010010101010101010100000000000000001011101110111011000000000000000001000100010001000000000000000000";
--X66Y57, nonlinear_LMDPL
constant Tile_X66Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000001011101110111011";
--X67Y57, linear_LMDPL
constant Tile_X67Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101010101011010101000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000011001100110011000000000000000000";
--X68Y57, linear_LMDPL
constant Tile_X68Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000101010100000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X69Y57, nonlinear_LMDPL
constant Tile_X69Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X70Y57, linear_LMDPL
constant Tile_X70Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000001011101110111011";
--X71Y57, linear_LMDPL
constant Tile_X71Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000001000100010001010011001100110010000000000000000";
--X72Y57, nonlinear_LMDPL
constant Tile_X72Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000001010101000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X73Y57, linear_LMDPL
constant Tile_X73Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000011111111000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000000100010001000110101010101010100000000000000000";
--X74Y57, linear_LMDPL
constant Tile_X74Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X75Y57, nonlinear_LMDPL
constant Tile_X75Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000001011101110111011";
--X76Y57, linear_LMDPL
constant Tile_X76Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010000010001000100010000000000000000";
--X77Y57, linear_LMDPL
constant Tile_X77Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000010001000100010";
--X78Y57, ctrl_to_sec
constant Tile_X78Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y57, combined_WDDL
constant Tile_X79Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y57, combined_WDDL
constant Tile_X80Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y57, ctrl_IO
constant Tile_X81Y57_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y58, W_IO_custom
constant Tile_X0Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y58, linear_LMDPL
constant Tile_X1Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010101010101010100000000000000001011101110111011000000000000000010001000100010000000000000000000";
--X2Y58, linear_LMDPL
constant Tile_X2Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010110101010000000000000000000000000101010100000000000000000010101010101010100000000000000001001100110011001000000000000000000000000000000000000000000000000";
--X3Y58, nonlinear_LMDPL
constant Tile_X3Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000110111011101110100000000000000001110111011101110";
--X4Y58, linear_LMDPL
constant Tile_X4Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000010001000100010010111011101110110000000000000000";
--X5Y58, linear_LMDPL
constant Tile_X5Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000110011001100110000100010001000100000000000000000";
--X6Y58, nonlinear_LMDPL
constant Tile_X6Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000101010110101010111111110000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100010001000100010000000000000000000";
--X7Y58, linear_LMDPL
constant Tile_X7Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100010001000100001010101010101010000000000000000";
--X8Y58, linear_LMDPL
constant Tile_X8Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010";
--X9Y58, nonlinear_LMDPL
constant Tile_X9Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001110111011101110";
--X10Y58, linear_LMDPL
constant Tile_X10Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000101010101010101001110111011101110000000000000000";
--X11Y58, linear_LMDPL
constant Tile_X11Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101010001000100010000000000000000000";
--X12Y58, nonlinear_LMDPL
constant Tile_X12Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000101010100000000000000000000000000000000000000001111111100000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000010001000100010000000000000000";
--X13Y58, linear_LMDPL
constant Tile_X13Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000000000000010101010101010100000000000000000000000000000000000000000000000001000100010001000000000000000000";
--X14Y58, linear_LMDPL
constant Tile_X14Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000100010001000110101010000000001000100010001000000000000000000000000000000000001000100010001000";
--X15Y58, nonlinear_LMDPL
constant Tile_X15Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000101010100000000011111111000000001010101000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000101010101010101011001100110011000000000000000000";
--X16Y58, linear_LMDPL
constant Tile_X16Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000100010001000100000000000000000000110011001100110";
--X17Y58, linear_LMDPL
constant Tile_X17Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X18Y58, nonlinear_LMDPL
constant Tile_X18Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000110111011101110110101010101010100000000000000000";
--X19Y58, linear_LMDPL
constant Tile_X19Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X20Y58, linear_LMDPL
constant Tile_X20Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000101010110101010010101010101010100000000000000000010001000100010000000000000000000110011001100110000000000000000";
--X21Y58, nonlinear_LMDPL
constant Tile_X21Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101011010101000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000101010100000000000000001010101000000000000000000000000000000000010101010101010100000000101010101010101010101010000000000000000010111011101110110000000000000000";
--X22Y58, linear_LMDPL
constant Tile_X22Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000011001100110011000000000000000001010101010101010000000000000000";
--X23Y58, linear_LMDPL
constant Tile_X23Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000101010100000000101010101010101001010101000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X24Y58, nonlinear_LMDPL
constant Tile_X24Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000010001000100010000000000101010100000000000000000001000100010001011001100110011000000000000000000";
--X25Y58, linear_LMDPL
constant Tile_X25Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X26Y58, linear_LMDPL
constant Tile_X26Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000010101010010101011010101000000000010101010101010100000000000000000010001000100010000000000000000001000100010001000000000000000000";
--X27Y58, nonlinear_LMDPL
constant Tile_X27Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101011010101000000000000000000000000000000000111111111010101000000000010101010000000000000000000000000000000010101010000000000101010100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101110111011101100000000000000000000000000000000";
--X28Y58, linear_LMDPL
constant Tile_X28Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000000101010100000000000000000000000010101010101010100101010110101010010101010101010100000000000000000110011001100110000000000000000010111011101110110000000000000000";
--X29Y58, linear_LMDPL
constant Tile_X29Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010101010100000000010101010101010100000000000000000000000000000000010101010000000001010101000000000101010100101010100000000000000000000000010101010010001000100010000000000101010100000000000000000001100110011001111001100110011000000000000000000";
--X30Y58, nonlinear_LMDPL
constant Tile_X30Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010100000000000000000000000001010101000000000000000000000000000000000101010101111111110101010000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X31Y58, linear_LMDPL
constant Tile_X31Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000101010100000000000000001010101011111111010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X32Y58, linear_LMDPL
constant Tile_X32Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000010101010111111110000000000000000101010100000000000000000000000000000000010101010010101010101010100000000000000001111111111111111000000000000000000000000000000000000000000000000";
--X33Y58, nonlinear_LMDPL
constant Tile_X33Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010101010000000000000000011111111000000000000000010101010101010101010101001010101000000001010101000000000101010100000000000000000000100010001000100000000101010100011001100110011000000000000000000000000000000000100010001000100";
--X34Y58, linear_LMDPL
constant Tile_X34Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101001010101111111110000000000000000000000000000000010101010000000000000000011111111010101010101010100000000000000000101010101010101000000000000000001000100010001000000000000000000";
--X35Y58, linear_LMDPL
constant Tile_X35Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101010101010101010000000000000000001010101000000000000000010101010000000000000000000000000010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X36Y58, nonlinear_LMDPL
constant Tile_X36Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000010101010101010100000000101010100010001000100010000000000000000010101010101010100000000000000000";
--X37Y58, linear_LMDPL
constant Tile_X37Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000000000000000000";
--X38Y58, linear_LMDPL
constant Tile_X38Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101011111111110101010000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010000000001010101000000000010001000100010000000000101010100000000000000000010001000100010011011101110111010000000000000000";
--X39Y58, nonlinear_LMDPL
constant Tile_X39Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000101010100000000000000001010101000000000000000001111111100000000000000000000000000000000101010100000000000000000001100110011001100000000000000000100010001000100";
--X40Y58, linear_LMDPL
constant Tile_X40Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000001111111111111111000000000000000011011101110111010000000000000000";
--X41Y58, linear_LMDPL
constant Tile_X41Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000001010101000100010001000100000000101010101010101010101010000000000000000000000000000000001110111011101110";
--X42Y58, nonlinear_LMDPL
constant Tile_X42Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010101010100000000010101010010101010101010100000000000000000010001000100010000000000000000010001000100010000000000000000000";
--X43Y58, linear_LMDPL
constant Tile_X43Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X44Y58, linear_LMDPL
constant Tile_X44Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000010101010101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000010101010000000000000000010101010010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X45Y58, nonlinear_LMDPL
constant Tile_X45Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010";
--X46Y58, linear_LMDPL
constant Tile_X46Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000000010001000100010";
--X47Y58, linear_LMDPL
constant Tile_X47Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111110101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101100000000000000000101010101010101";
--X48Y58, nonlinear_LMDPL
constant Tile_X48Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010001000100010000000000000000000000000000000000";
--X49Y58, linear_LMDPL
constant Tile_X49Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010000000001010101000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000010001000100010";
--X50Y58, linear_LMDPL
constant Tile_X50Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000010101010101010100000000000000001010101010101010000000000000000000000000000000000000000000000000";
--X51Y58, nonlinear_LMDPL
constant Tile_X51Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111111010101000000000010001000100010000000000101010100000000000000000001100110011001110001000100010000000000000000000";
--X52Y58, linear_LMDPL
constant Tile_X52Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X53Y58, linear_LMDPL
constant Tile_X53Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000101010100000000000000000000000000000000000000000000000000011001100110011";
--X54Y58, nonlinear_LMDPL
constant Tile_X54Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010101010101010100000000000000001000100010001000000000000000000011001100110011000000000000000000";
--X55Y58, linear_LMDPL
constant Tile_X55Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000101010101010101000110011001100110000000000000000";
--X56Y58, linear_LMDPL
constant Tile_X56Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X57Y58, nonlinear_LMDPL
constant Tile_X57Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000101010100000000000000000000000001010101000000000000000001111111100000000000000000000000000000000000000000000000000000000000100010001000100000000000000000100010001000100";
--X58Y58, linear_LMDPL
constant Tile_X58Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100";
--X59Y58, linear_LMDPL
constant Tile_X59Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X60Y58, nonlinear_LMDPL
constant Tile_X60Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001100100000000000000000101010101010101";
--X61Y58, linear_LMDPL
constant Tile_X61Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000001111111100000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X62Y58, linear_LMDPL
constant Tile_X62Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000010101010010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X63Y58, nonlinear_LMDPL
constant Tile_X63Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000001000100010001";
--X64Y58, linear_LMDPL
constant Tile_X64Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000011001100110011000000000000000000000000000000000101010101010101";
--X65Y58, linear_LMDPL
constant Tile_X65Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000101010100000000000000000101010101010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X66Y58, nonlinear_LMDPL
constant Tile_X66Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100100010001000100000000000000000010111011101110110000000000000000";
--X67Y58, linear_LMDPL
constant Tile_X67Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X68Y58, linear_LMDPL
constant Tile_X68Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101111111110000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000000100010001000100000000000000001000100010001000";
--X69Y58, nonlinear_LMDPL
constant Tile_X69Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000010001000100010";
--X70Y58, linear_LMDPL
constant Tile_X70Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010101010101010100000000000000000";
--X71Y58, linear_LMDPL
constant Tile_X71Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001001100110011001000000000000000000000000000000000001000100010001";
--X72Y58, nonlinear_LMDPL
constant Tile_X72Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101011111111010101010101010100000000000000001001100110011001000000000000000000010001000100010000000000000000";
--X73Y58, linear_LMDPL
constant Tile_X73Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000001000100010001000000000000000000000000000000000001011101110111011";
--X74Y58, linear_LMDPL
constant Tile_X74Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000001010101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000011111111010001000100010000000000000000000000000000000000010001000100010010001000100010000000000000000000";
--X75Y58, nonlinear_LMDPL
constant Tile_X75Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000101010111111111000000000000000001010101000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000001000100010001011001100110011000000000000000000";
--X76Y58, linear_LMDPL
constant Tile_X76Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111100000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001101110111011101000000000000000000000000000000000101010101010101";
--X77Y58, linear_LMDPL
constant Tile_X77Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000100010001000100000000000000001110111011101110000000000000000000000000000000000010001000100010";
--X78Y58, ctrl_to_sec
constant Tile_X78Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y58, combined_WDDL
constant Tile_X79Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y58, combined_WDDL
constant Tile_X80Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y58, ctrl_IO
constant Tile_X81Y58_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y59, W_IO_custom
constant Tile_X0Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y59, linear_LMDPL
constant Tile_X1Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000010101010111111110000000000000000010101010101010100000000000000000101010101010101000000000000000000010001000100010000000000000000";
--X2Y59, linear_LMDPL
constant Tile_X2Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X3Y59, nonlinear_LMDPL
constant Tile_X3Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000101010101010101010101010000000000000000010011001100110010000000000000000";
--X4Y59, linear_LMDPL
constant Tile_X4Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000010101010101010100000000000000001010101010101010000000000000000010001000100010000000000000000000";
--X5Y59, linear_LMDPL
constant Tile_X5Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X6Y59, nonlinear_LMDPL
constant Tile_X6Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001000100010001000";
--X7Y59, linear_LMDPL
constant Tile_X7Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100";
--X8Y59, linear_LMDPL
constant Tile_X8Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X9Y59, nonlinear_LMDPL
constant Tile_X9Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000001011101110111011";
--X10Y59, linear_LMDPL
constant Tile_X10Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000001010101000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X11Y59, linear_LMDPL
constant Tile_X11Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000100110011001100101110111011101110000000000000000";
--X12Y59, nonlinear_LMDPL
constant Tile_X12Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000000010001000100010000000000000000";
--X13Y59, linear_LMDPL
constant Tile_X13Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000101110111011101111001100110011000000000000000000";
--X14Y59, linear_LMDPL
constant Tile_X14Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000101010101010101000000000000000011011101110111010000000000000000";
--X15Y59, nonlinear_LMDPL
constant Tile_X15Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010011001100110010000000000000000";
--X16Y59, linear_LMDPL
constant Tile_X16Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000001010101000000000010101010000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100101010101010101000000000000000000100010001000100000000000000000";
--X17Y59, linear_LMDPL
constant Tile_X17Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X18Y59, nonlinear_LMDPL
constant Tile_X18Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010011001100110010000000000000000";
--X19Y59, linear_LMDPL
constant Tile_X19Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X20Y59, linear_LMDPL
constant Tile_X20Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000001000100010001000";
--X21Y59, nonlinear_LMDPL
constant Tile_X21Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X22Y59, linear_LMDPL
constant Tile_X22Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000010101011010101010101010000000000000000000000000000000001000100010001000";
--X23Y59, linear_LMDPL
constant Tile_X23Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000001010101000000000000000000000000101010100000000000000000101010100000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000010001000100010000000000000000000";
--X24Y59, nonlinear_LMDPL
constant Tile_X24Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000010101010000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100000000000000000000000000000000010111011101110110000000000000000";
--X25Y59, linear_LMDPL
constant Tile_X25Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101010100000000000000000000000000000000000000000000000011111111010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X26Y59, linear_LMDPL
constant Tile_X26Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000101010100000000000000000010101010101010100000000000000001011101110111011000000000000000011001100110011000000000000000000";
--X27Y59, nonlinear_LMDPL
constant Tile_X27Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010000000000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000010101010000000001010101000000000000000000000000000000000000000000101010100000000010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X28Y59, linear_LMDPL
constant Tile_X28Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000010101010101010100000000000000000101010100000000000000000000000001010101000000000000000000000000000000000111111111010101000000000000100010001000100000000000000001010101010101010000000000000000000000000000000000011001100110011";
--X29Y59, linear_LMDPL
constant Tile_X29Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101101010100000000000000000000000000000000011111111000000000000000001010101000000001010101000000000000000000000000010101010010001000100010000000000000000000000000000000000010001000100010000110011001100110000000000000000";
--X30Y59, nonlinear_LMDPL
constant Tile_X30Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000101010100000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010101010101010100000000000000000";
--X31Y59, linear_LMDPL
constant Tile_X31Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000001111111100000000000000000101010100000000000000000000000000000000000000001010101000000000010101010101010100000000000000000011001100110011000000000000000000100010001000100000000000000000";
--X32Y59, linear_LMDPL
constant Tile_X32Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000001010101000000000101010100000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000101010100000000000100010001000100000000000000000000000000000000000000000000000000000000000000001011101110111011";
--X33Y59, nonlinear_LMDPL
constant Tile_X33Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101000000000000000000000000000000000111111110000000001010101000000000000000000000000000000000000000001010101000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010101000100010001000000000000000000011001100110011000000000000000000";
--X34Y59, linear_LMDPL
constant Tile_X34Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010101010101010100000000000000000";
--X35Y59, linear_LMDPL
constant Tile_X35Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001000100010001000000000000000000000100010001000100000000000000000";
--X36Y59, nonlinear_LMDPL
constant Tile_X36Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101000000000000100010001000100000000101010100010001000100010000000000000000000000000000000000100010001000100";
--X37Y59, linear_LMDPL
constant Tile_X37Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010001000100010000000000000000000";
--X38Y59, linear_LMDPL
constant Tile_X38Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111101010100000000001010101000000000000000000000000000000000000000011111111000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X39Y59, nonlinear_LMDPL
constant Tile_X39Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X40Y59, linear_LMDPL
constant Tile_X40Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000001010101010101010000000000000000010111011101110110000000000000000";
--X41Y59, linear_LMDPL
constant Tile_X41Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000010101010010101010101010100000000101010101000100010001000000000000000000010101010101010100000000000000000";
--X42Y59, nonlinear_LMDPL
constant Tile_X42Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101010101010100000000101010101010101010101010000000000000000011001100110011000000000000000000";
--X43Y59, linear_LMDPL
constant Tile_X43Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000001000100010001010001000100010000000000000000000";
--X44Y59, linear_LMDPL
constant Tile_X44Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010111111110000000000000000000000000000000000000000000000001111111100000000000100010001000100000000000000001010101010101010000000000000000000000000000000000100010001000100";
--X45Y59, nonlinear_LMDPL
constant Tile_X45Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000001010101010101010";
--X46Y59, linear_LMDPL
constant Tile_X46Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000001010101010101010";
--X47Y59, linear_LMDPL
constant Tile_X47Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000110011001100110000000000000000";
--X48Y59, nonlinear_LMDPL
constant Tile_X48Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000110011001100110";
--X49Y59, linear_LMDPL
constant Tile_X49Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000010001000100010000000000000000000000000000000000110111011101110110111011101110110000000000000000";
--X50Y59, linear_LMDPL
constant Tile_X50Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010101010100000000000000000011001100110011000000000000000011001100110011000000000000000000";
--X51Y59, nonlinear_LMDPL
constant Tile_X51Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010001000100010000000000101010100000000000000000110111011101110110111011101110110000000000000000";
--X52Y59, linear_LMDPL
constant Tile_X52Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000100010001000100000000010101010010001000100010000000000000000000000000000000000100010001000100";
--X53Y59, linear_LMDPL
constant Tile_X53Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010001000100010000000000000000000000000000000000111011101110111011001100110011000000000000000000";
--X54Y59, nonlinear_LMDPL
constant Tile_X54Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100110000000000000000001001100110011001";
--X55Y59, linear_LMDPL
constant Tile_X55Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101010100000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000000100010001000100000000000000000";
--X56Y59, linear_LMDPL
constant Tile_X56Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010001000100010000000000000000000000000000000000110011001100110010101010101010100000000000000000";
--X57Y59, nonlinear_LMDPL
constant Tile_X57Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000111111110000000000000000000000000000000000000000000000000000000000000000000100010001000100000000101010101100110011001100000000000000000000000000000000001000100010001000";
--X58Y59, linear_LMDPL
constant Tile_X58Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000011001100110011";
--X59Y59, linear_LMDPL
constant Tile_X59Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001101110111011101000000000000000011111111111111110000000000000000";
--X60Y59, nonlinear_LMDPL
constant Tile_X60Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X61Y59, linear_LMDPL
constant Tile_X61Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000010011001100110010000000000000000";
--X62Y59, linear_LMDPL
constant Tile_X62Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100101010100000000010001000100010000000000000000000000000000000000011101110111011100110011001100110000000000000000";
--X63Y59, nonlinear_LMDPL
constant Tile_X63Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000001000100010001000000000000000000100010001000100";
--X64Y59, linear_LMDPL
constant Tile_X64Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011001100110011000100010001000100000000000000000";
--X65Y59, linear_LMDPL
constant Tile_X65Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000101010111111111000000000101010100000000000000000000000000000000000000001010101000000000101010100000000000000000000000001111111100000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000001000100010001000000000000000000011001100110011";
--X66Y59, nonlinear_LMDPL
constant Tile_X66Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000011111111000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000100010001000100000000000000001001100110011001000000000000000000000000000000000010001000100010";
--X67Y59, linear_LMDPL
constant Tile_X67Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000010101011010101000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011";
--X68Y59, linear_LMDPL
constant Tile_X68Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000101010100000000000000000101010100000000000000000111111111111111100000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110001000100010000000000000000000";
--X69Y59, nonlinear_LMDPL
constant Tile_X69Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000001100110011001100000000000000000001000100010001";
--X70Y59, linear_LMDPL
constant Tile_X70Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000101010101010101";
--X71Y59, linear_LMDPL
constant Tile_X71Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X72Y59, nonlinear_LMDPL
constant Tile_X72Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010101010101010100000000000000000";
--X73Y59, linear_LMDPL
constant Tile_X73Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000001010101000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000010001000100010000000000000000001010101010101010";
--X74Y59, linear_LMDPL
constant Tile_X74Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010010101010000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000110111011101110100000000000000000011001100110011";
--X75Y59, nonlinear_LMDPL
constant Tile_X75Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000010101010101010100000000000000000101010101010101000000000000000010001000100010000000000000000000";
--X76Y59, linear_LMDPL
constant Tile_X76Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000001111111100000000000000000000000010101010000000000000000000000000000000000000000000000000001000100010001000000000000000000000000000000000";
--X77Y59, linear_LMDPL
constant Tile_X77Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000110011001100110000000000000000010101010101010100000000000000000";
--X78Y59, ctrl_to_sec
constant Tile_X78Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y59, combined_WDDL
constant Tile_X79Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y59, combined_WDDL
constant Tile_X80Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y59, ctrl_IO
constant Tile_X81Y59_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X0Y60, W_IO_custom
constant Tile_X0Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X1Y60, linear_LMDPL
constant Tile_X1Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010001000100010000000000000000000";
--X2Y60, linear_LMDPL
constant Tile_X2Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000000000000000000000110011001100110000000000000000";
--X3Y60, nonlinear_LMDPL
constant Tile_X3Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X4Y60, linear_LMDPL
constant Tile_X4Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001101110111011101";
--X5Y60, linear_LMDPL
constant Tile_X5Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X6Y60, nonlinear_LMDPL
constant Tile_X6Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000010101010101010100000000000000000";
--X7Y60, linear_LMDPL
constant Tile_X7Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000001000100010001000000000000000000110011001100110000000000000000";
--X8Y60, linear_LMDPL
constant Tile_X8Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000011101110111011111001100110011000000000000000000";
--X9Y60, nonlinear_LMDPL
constant Tile_X9Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X10Y60, linear_LMDPL
constant Tile_X10Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001001100110011001000000000000000010111011101110110000000000000000";
--X11Y60, linear_LMDPL
constant Tile_X11Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010010011001100110010000000000000000";
--X12Y60, nonlinear_LMDPL
constant Tile_X12Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X13Y60, linear_LMDPL
constant Tile_X13Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000001010101010101010000000000000000000000000010001000100010000000000000000000000000000000000000000000000000001110111011101110000000000000000";
--X14Y60, linear_LMDPL
constant Tile_X14Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000010101010000000000000000000000000010101010101010100000000000000001100110011001100000000000000000001010101010101010000000000000000";
--X15Y60, nonlinear_LMDPL
constant Tile_X15Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000001000100010001000010001000100010000000000000000";
--X16Y60, linear_LMDPL
constant Tile_X16Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000101010101010101000000000000000000000000000000000010101010101010100000000000000000000000000000000000000000000000011011101110111010000000000000000";
--X17Y60, linear_LMDPL
constant Tile_X17Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X18Y60, nonlinear_LMDPL
constant Tile_X18Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X19Y60, linear_LMDPL
constant Tile_X19Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X20Y60, linear_LMDPL
constant Tile_X20Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X21Y60, nonlinear_LMDPL
constant Tile_X21Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X22Y60, linear_LMDPL
constant Tile_X22Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000001110111011101110";
--X23Y60, linear_LMDPL
constant Tile_X23Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001010101000000000000000000000000010101010101010100000000000000000010001000100010000000000000000001010101010101010000000000000000";
--X24Y60, nonlinear_LMDPL
constant Tile_X24Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011101110111011100000000000000000";
--X25Y60, linear_LMDPL
constant Tile_X25Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000101010100000000000000000000000001111111100000000000000001010101001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000110011001100110000000000000000000110011001100110000000000000000";
--X26Y60, linear_LMDPL
constant Tile_X26Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000100010001000100000000000000000011001100110011000000000000000000";
--X27Y60, nonlinear_LMDPL
constant Tile_X27Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000001010101000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000000000000000000000000000000000";
--X28Y60, linear_LMDPL
constant Tile_X28Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010101010000000000000000001010101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X29Y60, linear_LMDPL
constant Tile_X29Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000111111110000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010101010101010101010101010000000000000000000000000000000000000000000000000";
--X30Y60, nonlinear_LMDPL
constant Tile_X30Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X31Y60, linear_LMDPL
constant Tile_X31Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000101010101111111100000000000000000000000000000000000000000000000001010101000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000011001100110011000000000000000010111011101110110000000000000000";
--X32Y60, linear_LMDPL
constant Tile_X32Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000000000000000000000000000000000001010101010101010000000000000000";
--X33Y60, nonlinear_LMDPL
constant Tile_X33Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010100010001000100010000000000000000001110111011101110000000000000000";
--X34Y60, linear_LMDPL
constant Tile_X34Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000010001000100010000000000000000011011101110111010000000000000000";
--X35Y60, linear_LMDPL
constant Tile_X35Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000010101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101000000000000000000000000000000001101110111011101";
--X36Y60, nonlinear_LMDPL
constant Tile_X36Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010100101010101010101000000000000000010111011101110110000000000000000";
--X37Y60, linear_LMDPL
constant Tile_X37Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000";
--X38Y60, linear_LMDPL
constant Tile_X38Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X39Y60, nonlinear_LMDPL
constant Tile_X39Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X40Y60, linear_LMDPL
constant Tile_X40Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010111011101110110000000000000000";
--X41Y60, linear_LMDPL
constant Tile_X41Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000010101010101010100000000101010100011001100110011000000000000000010101010101010100000000000000000";
--X42Y60, nonlinear_LMDPL
constant Tile_X42Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X43Y60, linear_LMDPL
constant Tile_X43Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001111001100110011000000000000000000";
--X44Y60, linear_LMDPL
constant Tile_X44Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000010001000100010000000000000000000000000000000000";
--X45Y60, nonlinear_LMDPL
constant Tile_X45Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X46Y60, linear_LMDPL
constant Tile_X46Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X47Y60, linear_LMDPL
constant Tile_X47Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000010001000100010";
--X48Y60, nonlinear_LMDPL
constant Tile_X48Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X49Y60, linear_LMDPL
constant Tile_X49Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001000100010001000000000000000000010111011101110110000000000000000";
--X50Y60, linear_LMDPL
constant Tile_X50Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000010001000100010000000000000000000000000000000000010001000100010011001100110011000000000000000000";
--X51Y60, nonlinear_LMDPL
constant Tile_X51Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000";
--X52Y60, linear_LMDPL
constant Tile_X52Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000100010001000100";
--X53Y60, linear_LMDPL
constant Tile_X53Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000101010100000000000000000000000000000000011001100110011000000000000000000";
--X54Y60, nonlinear_LMDPL
constant Tile_X54Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010111011101110110000000000000000";
--X55Y60, linear_LMDPL
constant Tile_X55Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X56Y60, linear_LMDPL
constant Tile_X56Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X57Y60, nonlinear_LMDPL
constant Tile_X57Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000100010001000100";
--X58Y60, linear_LMDPL
constant Tile_X58Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110011";
--X59Y60, linear_LMDPL
constant Tile_X59Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X60Y60, nonlinear_LMDPL
constant Tile_X60Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X61Y60, linear_LMDPL
constant Tile_X61Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010110101010000000000010001000100010000000000000000010001000100010000000000000000000";
--X62Y60, linear_LMDPL
constant Tile_X62Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001100110011001100000000000000000010111011101110110000000000000000";
--X63Y60, nonlinear_LMDPL
constant Tile_X63Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X64Y60, linear_LMDPL
constant Tile_X64Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000000000000000000";
--X65Y60, linear_LMDPL
constant Tile_X65Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001100110011001100110011001100110000000000000000";
--X66Y60, nonlinear_LMDPL
constant Tile_X66Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000101010100010001000100010000000000000000001000100010001000000000000000000";
--X67Y60, linear_LMDPL
constant Tile_X67Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001001100110011001000000000000000010101010101010100000000000000000";
--X68Y60, linear_LMDPL
constant Tile_X68Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000010101010000000000000000101010100000000010101010000000000000000000000000000100010001000100000000000000001000100010001000000000000000000000000000000000000010001000100010";
--X69Y60, nonlinear_LMDPL
constant Tile_X69Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010001000100010000000000000000000000000000000000000100010001000110111011101110110000000000000000";
--X70Y60, linear_LMDPL
constant Tile_X70Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000100000000000000001101110111011101";
--X71Y60, linear_LMDPL
constant Tile_X71Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011001100000000000000000010001000100010";
--X72Y60, nonlinear_LMDPL
constant Tile_X72Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X73Y60, linear_LMDPL
constant Tile_X73Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000001011101110111011000000000000000000110011001100110000000000000000";
--X74Y60, linear_LMDPL
constant Tile_X74Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000000000000000000000010101010101010100000000000000001100110011001100000000000000000000000000000000000000000000000000";
--X75Y60, nonlinear_LMDPL
constant Tile_X75Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010100000000000000000100010001000100000000000000000010111011101110110000000000000000";
--X76Y60, linear_LMDPL
constant Tile_X76Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100010000000000000000000000000000000000001000100010001010101010101010100000000000000000";
--X77Y60, linear_LMDPL
constant Tile_X77Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X78Y60, ctrl_to_sec
constant Tile_X78Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X79Y60, combined_WDDL
constant Tile_X79Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X80Y60, combined_WDDL
constant Tile_X80Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--X81Y60, ctrl_IO
constant Tile_X81Y60_Emulate_Bitstream : std_logic_vector(640-1 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
end package emulate_bitstream;
