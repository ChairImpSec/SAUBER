/* modified netlist. Source: module present in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/11-PRESENT80_nibble_serial_encryption_PortParallel/4-AGEMA/present.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module present_SAUBER_Pipeline_d1 (data_in_s0_t, key_s0_t, reset_t, data_in_s0_f, data_in_s1_t, data_in_s1_f, key_s0_f, key_s1_t, key_s1_f, reset_f, data_out_s0_t, done_t, data_out_s0_f, data_out_s1_t, data_out_s1_f, done_f);
    input [63:0] data_in_s0_t ;
    input [79:0] key_s0_t ;
    input reset_t ;
    input [63:0] data_in_s0_f ;
    input [63:0] data_in_s1_t ;
    input [63:0] data_in_s1_f ;
    input [79:0] key_s0_f ;
    input [79:0] key_s1_t ;
    input [79:0] key_s1_f ;
    input reset_f ;
    output [63:0] data_out_s0_t ;
    output done_t ;
    output [63:0] data_out_s0_f ;
    output [63:0] data_out_s1_t ;
    output [63:0] data_out_s1_f ;
    output done_f ;
    wire selSbox ;
    wire intDone ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n5 ;
    wire fsm_n4 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_n16 ;
    wire fsm_ps_state_0_ ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n4 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n2 ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y ;
    wire stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_0_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_0_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_1_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_1_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_2_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_2_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_3_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_3_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_4_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_4_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_5_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_5_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_6_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_6_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_7_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_7_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_8_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_8_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_9_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_9_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_10_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_10_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_11_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_11_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_12_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_12_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_13_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_13_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_14_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_14_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_15_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_15_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_16_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_16_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_17_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_17_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_18_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_18_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_19_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_19_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_20_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_20_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_21_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_21_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_22_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_22_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_23_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_23_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_24_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_24_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_25_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_25_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_26_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_26_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_27_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_27_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_28_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_28_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_29_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_29_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_30_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_30_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_31_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_31_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_32_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_32_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_33_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_33_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_34_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_34_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_35_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_35_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_36_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_36_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_37_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_37_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_38_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_38_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_39_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_39_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_40_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_40_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_41_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_41_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_42_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_42_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_43_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_43_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_44_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_44_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_45_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_45_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_46_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_46_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_47_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_47_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_48_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_48_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_49_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_49_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_50_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_50_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_51_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_51_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_52_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_52_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_53_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_53_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_54_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_54_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_55_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_55_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_56_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_56_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_57_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_57_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_58_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_58_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_59_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_59_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_60_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_60_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_61_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_61_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_62_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_62_U1_X ;
    wire stateFF_MUX_inputPar_mux_inst_63_U1_Y ;
    wire stateFF_MUX_inputPar_mux_inst_63_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y ;
    wire keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_0_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_0_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_1_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_1_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_2_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_2_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_3_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_3_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_4_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_4_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_5_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_5_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_6_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_6_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_7_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_7_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_8_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_8_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_9_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_9_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_10_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_10_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_11_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_11_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_12_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_12_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_13_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_13_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_14_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_14_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_15_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_15_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_16_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_16_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_17_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_17_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_18_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_18_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_19_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_19_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_20_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_20_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_21_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_21_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_22_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_22_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_23_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_23_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_24_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_24_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_25_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_25_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_26_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_26_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_27_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_27_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_28_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_28_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_29_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_29_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_30_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_30_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_31_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_31_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_32_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_32_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_33_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_33_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_34_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_34_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_35_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_35_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_36_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_36_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_37_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_37_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_38_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_38_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_39_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_39_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_40_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_40_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_41_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_41_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_42_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_42_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_43_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_43_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_44_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_44_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_45_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_45_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_46_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_46_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_47_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_47_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_48_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_48_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_49_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_49_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_50_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_50_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_51_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_51_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_52_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_52_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_53_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_53_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_54_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_54_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_55_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_55_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_56_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_56_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_57_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_57_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_58_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_58_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_59_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_59_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_60_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_60_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_61_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_61_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_62_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_62_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_63_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_63_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_64_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_64_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_65_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_65_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_66_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_66_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_67_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_67_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_68_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_68_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_69_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_69_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_70_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_70_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_71_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_71_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_72_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_72_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_73_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_73_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_74_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_74_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_75_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_75_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_76_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_76_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_77_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_77_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_78_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_78_U1_X ;
    wire keyFF_MUX_inputPar_mux_inst_79_U1_Y ;
    wire keyFF_MUX_inputPar_mux_inst_79_U1_X ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire MUX_sboxin_mux_inst_0_U1_Y ;
    wire MUX_sboxin_mux_inst_0_U1_X ;
    wire MUX_sboxin_mux_inst_1_U1_Y ;
    wire MUX_sboxin_mux_inst_1_U1_X ;
    wire MUX_sboxin_mux_inst_2_U1_Y ;
    wire MUX_sboxin_mux_inst_2_U1_X ;
    wire MUX_sboxin_mux_inst_3_U1_Y ;
    wire MUX_sboxin_mux_inst_3_U1_X ;
    wire MUX_serialIn_mux_inst_0_U1_Y ;
    wire MUX_serialIn_mux_inst_0_U1_X ;
    wire MUX_serialIn_mux_inst_1_U1_Y ;
    wire MUX_serialIn_mux_inst_1_U1_X ;
    wire MUX_serialIn_mux_inst_2_U1_Y ;
    wire MUX_serialIn_mux_inst_2_U1_X ;
    wire MUX_serialIn_mux_inst_3_U1_Y ;
    wire MUX_serialIn_mux_inst_3_U1_X ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2136 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2140 ;
    wire new_AGEMA_signal_2144 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2334 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2482 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2488 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2500 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2506 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2518 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2524 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2536 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2542 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2554 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2560 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2572 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2850 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2856 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2862 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2868 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2876 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2882 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2888 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2894 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2900 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2906 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2912 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2918 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U9 ( .A0_t (roundkey[1]), .A0_f (new_AGEMA_signal_1434), .A1_t (new_AGEMA_signal_1435), .A1_f (new_AGEMA_signal_1436), .B0_t (data_out_s0_t[61]), .B0_f (data_out_s0_f[61]), .B1_t (data_out_s1_t[61]), .B1_f (data_out_s1_f[61]), .Z0_t (stateXORroundkey[1]), .Z0_f (new_AGEMA_signal_1440), .Z1_t (new_AGEMA_signal_1441), .Z1_f (new_AGEMA_signal_1442) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U10 ( .A0_t (roundkey[2]), .A0_f (new_AGEMA_signal_1443), .A1_t (new_AGEMA_signal_1444), .A1_f (new_AGEMA_signal_1445), .B0_t (data_out_s0_t[62]), .B0_f (data_out_s0_f[62]), .B1_t (data_out_s1_t[62]), .B1_f (data_out_s1_f[62]), .Z0_t (stateXORroundkey[2]), .Z0_f (new_AGEMA_signal_1449), .Z1_t (new_AGEMA_signal_1450), .Z1_f (new_AGEMA_signal_1451) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U11 ( .A0_t (roundkey[0]), .A0_f (new_AGEMA_signal_1452), .A1_t (new_AGEMA_signal_1453), .A1_f (new_AGEMA_signal_1454), .B0_t (data_out_s0_t[60]), .B0_f (data_out_s0_f[60]), .B1_t (data_out_s1_t[60]), .B1_f (data_out_s1_f[60]), .Z0_t (stateXORroundkey[0]), .Z0_f (new_AGEMA_signal_1458), .Z1_t (new_AGEMA_signal_1459), .Z1_f (new_AGEMA_signal_1460) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) U12 ( .A0_t (roundkey[3]), .A0_f (new_AGEMA_signal_1461), .A1_t (new_AGEMA_signal_1462), .A1_f (new_AGEMA_signal_1463), .B0_t (data_out_s0_t[63]), .B0_f (data_out_s0_f[63]), .B1_t (data_out_s1_t[63]), .B1_f (data_out_s1_f[63]), .Z0_t (stateXORroundkey[3]), .Z0_f (new_AGEMA_signal_1467), .Z1_t (new_AGEMA_signal_1468), .Z1_f (new_AGEMA_signal_1469) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_U19 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (fsm_n14), .B0_f (new_AGEMA_signal_3613), .Z0_t (fsm_n16), .Z0_f (new_AGEMA_signal_1479) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U18 ( .A0_t (fsm_n16), .A0_f (new_AGEMA_signal_1479), .B0_t (fsm_n13), .B0_f (new_AGEMA_signal_3177), .Z0_t (fsm_n14), .Z0_f (new_AGEMA_signal_3613) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U17 ( .A0_t (fsm_n12), .A0_f (new_AGEMA_signal_2714), .B0_t (fsm_n11), .B0_f (new_AGEMA_signal_1472), .Z0_t (fsm_n13), .Z0_f (new_AGEMA_signal_3177) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U16 ( .A0_t (counter[3]), .A0_f (new_AGEMA_signal_1470), .B0_t (fsm_ps_state_0_), .B0_f (new_AGEMA_signal_1471), .Z0_t (fsm_n11), .Z0_f (new_AGEMA_signal_1472) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U15 ( .A0_t (fsm_n10), .A0_f (new_AGEMA_signal_1478), .B0_t (fsm_n9), .B0_f (new_AGEMA_signal_1475), .Z0_t (fsm_n12), .Z0_f (new_AGEMA_signal_2714) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U14 ( .A0_t (counter[4]), .A0_f (new_AGEMA_signal_1473), .B0_t (counter[0]), .B0_f (new_AGEMA_signal_1474), .Z0_t (fsm_n9), .Z0_f (new_AGEMA_signal_1475) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U13 ( .A0_t (counter[1]), .A0_f (new_AGEMA_signal_1476), .B0_t (counter[2]), .B0_f (new_AGEMA_signal_1477), .Z0_t (fsm_n10), .Z0_f (new_AGEMA_signal_1478) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U12 ( .A0_t (fsm_n16), .A0_f (new_AGEMA_signal_1479), .B0_t (fsm_ps_state_0_), .B0_f (new_AGEMA_signal_1471), .Z0_t (intDone), .Z0_f (new_AGEMA_signal_1480) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U11 ( .A0_t (fsm_n8), .A0_f (new_AGEMA_signal_3178), .B0_t (fsm_n16), .B0_f (new_AGEMA_signal_1479), .Z0_t (fsm_en_countRound), .Z0_f (new_AGEMA_signal_3614) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_U10 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (fsm_n7), .B0_f (new_AGEMA_signal_3615), .Z0_t (fsm_ps_state_0_), .Z0_f (new_AGEMA_signal_1471) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U9 ( .A0_t (fsm_n8), .A0_f (new_AGEMA_signal_3178), .B0_t (done_t), .B0_f (done_f), .Z0_t (fsm_n7), .Z0_f (new_AGEMA_signal_3615) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U8 ( .A0_t (fsm_countSerial[1]), .A0_f (new_AGEMA_signal_2718), .B0_t (fsm_n6), .B0_f (new_AGEMA_signal_2715), .Z0_t (fsm_n8), .Z0_f (new_AGEMA_signal_3178) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U7 ( .A0_t (fsm_n5), .A0_f (new_AGEMA_signal_1485), .B0_t (fsm_n4), .B0_f (new_AGEMA_signal_1483), .Z0_t (fsm_n6), .Z0_f (new_AGEMA_signal_2715) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U6 ( .A0_t (fsm_countSerial[3]), .A0_f (new_AGEMA_signal_1481), .B0_t (fsm_countSerial[2]), .B0_f (new_AGEMA_signal_1482), .Z0_t (fsm_n4), .Z0_f (new_AGEMA_signal_1483) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_U5 ( .A0_t (fsm_ps_state_0_), .A0_f (new_AGEMA_signal_1471), .B0_t (fsm_countSerial[0]), .B0_f (new_AGEMA_signal_1484), .Z0_t (fsm_n5), .Z0_f (new_AGEMA_signal_1485) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U4 ( .A0_t (fsm_ps_state_0_), .A0_f (new_AGEMA_signal_1471), .B0_t (fsm_n16), .B0_f (new_AGEMA_signal_1479), .Z0_t (done_t), .Z0_f (done_f) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U2 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (selSbox), .B0_f (new_AGEMA_signal_1487), .Z0_t (fsm_rst_countSerial), .Z0_f (new_AGEMA_signal_2717) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_U1 ( .A0_t (fsm_ps_state_0_), .A0_f (new_AGEMA_signal_1471), .B0_t (fsm_n16), .B0_f (new_AGEMA_signal_1479), .Z0_t (selSbox), .Z0_f (new_AGEMA_signal_1487) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U15 ( .A0_t (fsm_cnt_rnd_n12), .A0_f (new_AGEMA_signal_4494), .B0_t (reset_t), .B0_f (reset_f), .Z0_t (counter[2]), .Z0_f (new_AGEMA_signal_1477) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U14 ( .A0_t (fsm_cnt_rnd_n10), .A0_f (new_AGEMA_signal_4463), .B0_t (counter[2]), .B0_f (new_AGEMA_signal_1477), .Z0_t (fsm_cnt_rnd_n12), .Z0_f (new_AGEMA_signal_4494) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U13 ( .A0_t (fsm_cnt_rnd_n9), .A0_f (new_AGEMA_signal_4037), .B0_t (reset_t), .B0_f (reset_f), .Z0_t (counter[0]), .Z0_f (new_AGEMA_signal_1474) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U12 ( .A0_t (counter[0]), .A0_f (new_AGEMA_signal_1474), .B0_t (fsm_en_countRound), .B0_f (new_AGEMA_signal_3614), .Z0_t (fsm_cnt_rnd_n9), .Z0_f (new_AGEMA_signal_4037) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U11 ( .A0_t (fsm_cnt_rnd_n8), .A0_f (new_AGEMA_signal_4525), .B0_t (reset_t), .B0_f (reset_f), .Z0_t (counter[4]), .Z0_f (new_AGEMA_signal_1473) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U10 ( .A0_t (counter[4]), .A0_f (new_AGEMA_signal_1473), .B0_t (fsm_cnt_rnd_n7), .B0_f (new_AGEMA_signal_4511), .Z0_t (fsm_cnt_rnd_n8), .Z0_f (new_AGEMA_signal_4525) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U9 ( .A0_t (counter[3]), .A0_f (new_AGEMA_signal_1470), .B0_t (fsm_cnt_rnd_n6), .B0_f (new_AGEMA_signal_4495), .Z0_t (fsm_cnt_rnd_n7), .Z0_f (new_AGEMA_signal_4511) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U8 ( .A0_t (reset_t), .A0_f (reset_f), .B0_t (fsm_cnt_rnd_n5), .B0_f (new_AGEMA_signal_4462), .Z0_t (counter[1]), .Z0_f (new_AGEMA_signal_1476) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U7 ( .A0_t (counter[1]), .A0_f (new_AGEMA_signal_1476), .B0_t (fsm_cnt_rnd_n4), .B0_f (new_AGEMA_signal_4038), .Z0_t (fsm_cnt_rnd_n5), .Z0_f (new_AGEMA_signal_4462) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_rnd_U6 ( .A0_t (fsm_cnt_rnd_n3), .A0_f (new_AGEMA_signal_4512), .B0_t (reset_t), .B0_f (reset_f), .Z0_t (counter[3]), .Z0_f (new_AGEMA_signal_1470) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_rnd_U4 ( .A0_t (fsm_cnt_rnd_n6), .A0_f (new_AGEMA_signal_4495), .B0_t (counter[3]), .B0_f (new_AGEMA_signal_1470), .Z0_t (fsm_cnt_rnd_n3), .Z0_f (new_AGEMA_signal_4512) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U3 ( .A0_t (fsm_cnt_rnd_n10), .A0_f (new_AGEMA_signal_4463), .B0_t (counter[2]), .B0_f (new_AGEMA_signal_1477), .Z0_t (fsm_cnt_rnd_n6), .Z0_f (new_AGEMA_signal_4495) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U2 ( .A0_t (counter[1]), .A0_f (new_AGEMA_signal_1476), .B0_t (fsm_cnt_rnd_n4), .B0_f (new_AGEMA_signal_4038), .Z0_t (fsm_cnt_rnd_n10), .Z0_f (new_AGEMA_signal_4463) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_rnd_U1 ( .A0_t (counter[0]), .A0_f (new_AGEMA_signal_1474), .B0_t (fsm_en_countRound), .B0_f (new_AGEMA_signal_3614), .Z0_t (fsm_cnt_rnd_n4), .Z0_f (new_AGEMA_signal_4038) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U12 ( .A0_t (fsm_cnt_ser_n9), .A0_f (new_AGEMA_signal_1488), .B0_t (fsm_rst_countSerial), .B0_f (new_AGEMA_signal_2717), .Z0_t (fsm_countSerial[0]), .Z0_f (new_AGEMA_signal_1484) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U11 ( .A0_t (fsm_ps_state_0_), .A0_f (new_AGEMA_signal_1471), .B0_t (fsm_countSerial[0]), .B0_f (new_AGEMA_signal_1484), .Z0_t (fsm_cnt_ser_n9), .Z0_f (new_AGEMA_signal_1488) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U10 ( .A0_t (fsm_cnt_ser_n7), .A0_f (new_AGEMA_signal_2719), .B0_t (fsm_rst_countSerial), .B0_f (new_AGEMA_signal_2717), .Z0_t (fsm_countSerial[1]), .Z0_f (new_AGEMA_signal_2718) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U9 ( .A0_t (fsm_cnt_ser_n6), .A0_f (new_AGEMA_signal_1489), .B0_t (fsm_countSerial[1]), .B0_f (new_AGEMA_signal_2718), .Z0_t (fsm_cnt_ser_n7), .Z0_f (new_AGEMA_signal_2719) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U8 ( .A0_t (fsm_cnt_ser_n5), .A0_f (new_AGEMA_signal_3616), .B0_t (fsm_rst_countSerial), .B0_f (new_AGEMA_signal_2717), .Z0_t (fsm_countSerial[3]), .Z0_f (new_AGEMA_signal_1481) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U7 ( .A0_t (fsm_countSerial[3]), .A0_f (new_AGEMA_signal_1481), .B0_t (fsm_cnt_ser_n4), .B0_f (new_AGEMA_signal_3179), .Z0_t (fsm_cnt_ser_n5), .Z0_f (new_AGEMA_signal_3616) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U6 ( .A0_t (fsm_countSerial[2]), .A0_f (new_AGEMA_signal_1482), .B0_t (fsm_cnt_ser_n3), .B0_f (new_AGEMA_signal_2720), .Z0_t (fsm_cnt_ser_n4), .Z0_f (new_AGEMA_signal_3179) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b1)) fsm_cnt_ser_U5 ( .A0_t (fsm_cnt_ser_n2), .A0_f (new_AGEMA_signal_3180), .B0_t (fsm_rst_countSerial), .B0_f (new_AGEMA_signal_2717), .Z0_t (fsm_countSerial[2]), .Z0_f (new_AGEMA_signal_1482) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b0)) fsm_cnt_ser_U3 ( .A0_t (fsm_cnt_ser_n3), .A0_f (new_AGEMA_signal_2720), .B0_t (fsm_countSerial[2]), .B0_f (new_AGEMA_signal_1482), .Z0_t (fsm_cnt_ser_n2), .Z0_f (new_AGEMA_signal_3180) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U2 ( .A0_t (fsm_cnt_ser_n6), .A0_f (new_AGEMA_signal_1489), .B0_t (fsm_countSerial[1]), .B0_f (new_AGEMA_signal_2718), .Z0_t (fsm_cnt_ser_n3), .Z0_f (new_AGEMA_signal_2720) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) fsm_cnt_ser_U1 ( .A0_t (fsm_ps_state_0_), .A0_f (new_AGEMA_signal_1471), .B0_t (fsm_countSerial[0]), .B0_f (new_AGEMA_signal_1484), .Z0_t (fsm_cnt_ser_n6), .Z0_f (new_AGEMA_signal_1489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (serialIn[0]), .A0_f (new_AGEMA_signal_4535), .A1_t (new_AGEMA_signal_4536), .A1_f (new_AGEMA_signal_4537), .B0_t (stateFF_inputPar[0]), .B0_f (new_AGEMA_signal_3181), .B1_t (new_AGEMA_signal_3182), .B1_f (new_AGEMA_signal_3183), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_4538), .Z1_t (new_AGEMA_signal_4539), .Z1_f (new_AGEMA_signal_4540) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_4538), .B1_t (new_AGEMA_signal_4539), .B1_f (new_AGEMA_signal_4540), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4553), .Z1_t (new_AGEMA_signal_4554), .Z1_f (new_AGEMA_signal_4555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4553), .A1_t (new_AGEMA_signal_4554), .A1_f (new_AGEMA_signal_4555), .B0_t (serialIn[0]), .B0_f (new_AGEMA_signal_4535), .B1_t (new_AGEMA_signal_4536), .B1_f (new_AGEMA_signal_4537), .Z0_t (data_out_s0_t[0]), .Z0_f (data_out_s0_f[0]), .Z1_t (data_out_s1_t[0]), .Z1_f (data_out_s1_f[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (serialIn[1]), .A0_f (new_AGEMA_signal_4610), .A1_t (new_AGEMA_signal_4611), .A1_f (new_AGEMA_signal_4612), .B0_t (stateFF_inputPar[1]), .B0_f (new_AGEMA_signal_3184), .B1_t (new_AGEMA_signal_3185), .B1_f (new_AGEMA_signal_3186), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4619), .Z1_t (new_AGEMA_signal_4620), .Z1_f (new_AGEMA_signal_4621) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4619), .B1_t (new_AGEMA_signal_4620), .B1_f (new_AGEMA_signal_4621), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4637), .Z1_t (new_AGEMA_signal_4638), .Z1_f (new_AGEMA_signal_4639) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4637), .A1_t (new_AGEMA_signal_4638), .A1_f (new_AGEMA_signal_4639), .B0_t (serialIn[1]), .B0_f (new_AGEMA_signal_4610), .B1_t (new_AGEMA_signal_4611), .B1_f (new_AGEMA_signal_4612), .Z0_t (data_out_s0_t[1]), .Z0_f (data_out_s0_f[1]), .Z1_t (data_out_s1_t[1]), .Z1_f (data_out_s1_f[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (serialIn[2]), .A0_f (new_AGEMA_signal_4613), .A1_t (new_AGEMA_signal_4614), .A1_f (new_AGEMA_signal_4615), .B0_t (stateFF_inputPar[2]), .B0_f (new_AGEMA_signal_3187), .B1_t (new_AGEMA_signal_3188), .B1_f (new_AGEMA_signal_3189), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_4622), .Z1_t (new_AGEMA_signal_4623), .Z1_f (new_AGEMA_signal_4624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_4622), .B1_t (new_AGEMA_signal_4623), .B1_f (new_AGEMA_signal_4624), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4640), .Z1_t (new_AGEMA_signal_4641), .Z1_f (new_AGEMA_signal_4642) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4640), .A1_t (new_AGEMA_signal_4641), .A1_f (new_AGEMA_signal_4642), .B0_t (serialIn[2]), .B0_f (new_AGEMA_signal_4613), .B1_t (new_AGEMA_signal_4614), .B1_f (new_AGEMA_signal_4615), .Z0_t (data_out_s0_t[2]), .Z0_f (data_out_s0_f[2]), .Z1_t (data_out_s1_t[2]), .Z1_f (data_out_s1_f[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (serialIn[3]), .A0_f (new_AGEMA_signal_4634), .A1_t (new_AGEMA_signal_4635), .A1_f (new_AGEMA_signal_4636), .B0_t (stateFF_inputPar[3]), .B0_f (new_AGEMA_signal_3190), .B1_t (new_AGEMA_signal_3191), .B1_f (new_AGEMA_signal_3192), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4643), .Z1_t (new_AGEMA_signal_4644), .Z1_f (new_AGEMA_signal_4645) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4643), .B1_t (new_AGEMA_signal_4644), .B1_f (new_AGEMA_signal_4645), .Z0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4655), .Z1_t (new_AGEMA_signal_4656), .Z1_f (new_AGEMA_signal_4657) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4655), .A1_t (new_AGEMA_signal_4656), .A1_f (new_AGEMA_signal_4657), .B0_t (serialIn[3]), .B0_f (new_AGEMA_signal_4634), .B1_t (new_AGEMA_signal_4635), .B1_f (new_AGEMA_signal_4636), .Z0_t (data_out_s0_t[3]), .Z0_f (data_out_s0_f[3]), .Z1_t (data_out_s1_t[3]), .Z1_f (data_out_s1_f[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[0]), .A0_f (data_out_s0_f[0]), .A1_t (data_out_s1_t[0]), .A1_f (data_out_s1_f[0]), .B0_t (stateFF_inputPar[4]), .B0_f (new_AGEMA_signal_3193), .B1_t (new_AGEMA_signal_3194), .B1_f (new_AGEMA_signal_3195), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3617), .Z1_t (new_AGEMA_signal_3618), .Z1_f (new_AGEMA_signal_3619) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3617), .B1_t (new_AGEMA_signal_3618), .B1_f (new_AGEMA_signal_3619), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4039), .Z1_t (new_AGEMA_signal_4040), .Z1_f (new_AGEMA_signal_4041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4039), .A1_t (new_AGEMA_signal_4040), .A1_f (new_AGEMA_signal_4041), .B0_t (data_out_s0_t[0]), .B0_f (data_out_s0_f[0]), .B1_t (data_out_s1_t[0]), .B1_f (data_out_s1_f[0]), .Z0_t (data_out_s0_t[4]), .Z0_f (data_out_s0_f[4]), .Z1_t (data_out_s1_t[4]), .Z1_f (data_out_s1_f[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[1]), .A0_f (data_out_s0_f[1]), .A1_t (data_out_s1_t[1]), .A1_f (data_out_s1_f[1]), .B0_t (stateFF_inputPar[5]), .B0_f (new_AGEMA_signal_3196), .B1_t (new_AGEMA_signal_3197), .B1_f (new_AGEMA_signal_3198), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3620), .Z1_t (new_AGEMA_signal_3621), .Z1_f (new_AGEMA_signal_3622) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3620), .B1_t (new_AGEMA_signal_3621), .B1_f (new_AGEMA_signal_3622), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4042), .Z1_t (new_AGEMA_signal_4043), .Z1_f (new_AGEMA_signal_4044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4042), .A1_t (new_AGEMA_signal_4043), .A1_f (new_AGEMA_signal_4044), .B0_t (data_out_s0_t[1]), .B0_f (data_out_s0_f[1]), .B1_t (data_out_s1_t[1]), .B1_f (data_out_s1_f[1]), .Z0_t (data_out_s0_t[5]), .Z0_f (data_out_s0_f[5]), .Z1_t (data_out_s1_t[5]), .Z1_f (data_out_s1_f[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[2]), .A0_f (data_out_s0_f[2]), .A1_t (data_out_s1_t[2]), .A1_f (data_out_s1_f[2]), .B0_t (stateFF_inputPar[6]), .B0_f (new_AGEMA_signal_3199), .B1_t (new_AGEMA_signal_3200), .B1_f (new_AGEMA_signal_3201), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3623), .Z1_t (new_AGEMA_signal_3624), .Z1_f (new_AGEMA_signal_3625) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3623), .B1_t (new_AGEMA_signal_3624), .B1_f (new_AGEMA_signal_3625), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4045), .Z1_t (new_AGEMA_signal_4046), .Z1_f (new_AGEMA_signal_4047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4045), .A1_t (new_AGEMA_signal_4046), .A1_f (new_AGEMA_signal_4047), .B0_t (data_out_s0_t[2]), .B0_f (data_out_s0_f[2]), .B1_t (data_out_s1_t[2]), .B1_f (data_out_s1_f[2]), .Z0_t (data_out_s0_t[6]), .Z0_f (data_out_s0_f[6]), .Z1_t (data_out_s1_t[6]), .Z1_f (data_out_s1_f[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[3]), .A0_f (data_out_s0_f[3]), .A1_t (data_out_s1_t[3]), .A1_f (data_out_s1_f[3]), .B0_t (stateFF_inputPar[7]), .B0_f (new_AGEMA_signal_3202), .B1_t (new_AGEMA_signal_3203), .B1_f (new_AGEMA_signal_3204), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3626), .Z1_t (new_AGEMA_signal_3627), .Z1_f (new_AGEMA_signal_3628) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3626), .B1_t (new_AGEMA_signal_3627), .B1_f (new_AGEMA_signal_3628), .Z0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4048), .Z1_t (new_AGEMA_signal_4049), .Z1_f (new_AGEMA_signal_4050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4048), .A1_t (new_AGEMA_signal_4049), .A1_f (new_AGEMA_signal_4050), .B0_t (data_out_s0_t[3]), .B0_f (data_out_s0_f[3]), .B1_t (data_out_s1_t[3]), .B1_f (data_out_s1_f[3]), .Z0_t (data_out_s0_t[7]), .Z0_f (data_out_s0_f[7]), .Z1_t (data_out_s1_t[7]), .Z1_f (data_out_s1_f[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[4]), .A0_f (data_out_s0_f[4]), .A1_t (data_out_s1_t[4]), .A1_f (data_out_s1_f[4]), .B0_t (stateFF_inputPar[8]), .B0_f (new_AGEMA_signal_3205), .B1_t (new_AGEMA_signal_3206), .B1_f (new_AGEMA_signal_3207), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3629), .Z1_t (new_AGEMA_signal_3630), .Z1_f (new_AGEMA_signal_3631) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3629), .B1_t (new_AGEMA_signal_3630), .B1_f (new_AGEMA_signal_3631), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4051), .Z1_t (new_AGEMA_signal_4052), .Z1_f (new_AGEMA_signal_4053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4051), .A1_t (new_AGEMA_signal_4052), .A1_f (new_AGEMA_signal_4053), .B0_t (data_out_s0_t[4]), .B0_f (data_out_s0_f[4]), .B1_t (data_out_s1_t[4]), .B1_f (data_out_s1_f[4]), .Z0_t (data_out_s0_t[8]), .Z0_f (data_out_s0_f[8]), .Z1_t (data_out_s1_t[8]), .Z1_f (data_out_s1_f[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[5]), .A0_f (data_out_s0_f[5]), .A1_t (data_out_s1_t[5]), .A1_f (data_out_s1_f[5]), .B0_t (stateFF_inputPar[9]), .B0_f (new_AGEMA_signal_3208), .B1_t (new_AGEMA_signal_3209), .B1_f (new_AGEMA_signal_3210), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3632), .Z1_t (new_AGEMA_signal_3633), .Z1_f (new_AGEMA_signal_3634) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3632), .B1_t (new_AGEMA_signal_3633), .B1_f (new_AGEMA_signal_3634), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4054), .Z1_t (new_AGEMA_signal_4055), .Z1_f (new_AGEMA_signal_4056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4054), .A1_t (new_AGEMA_signal_4055), .A1_f (new_AGEMA_signal_4056), .B0_t (data_out_s0_t[5]), .B0_f (data_out_s0_f[5]), .B1_t (data_out_s1_t[5]), .B1_f (data_out_s1_f[5]), .Z0_t (data_out_s0_t[9]), .Z0_f (data_out_s0_f[9]), .Z1_t (data_out_s1_t[9]), .Z1_f (data_out_s1_f[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[6]), .A0_f (data_out_s0_f[6]), .A1_t (data_out_s1_t[6]), .A1_f (data_out_s1_f[6]), .B0_t (stateFF_inputPar[10]), .B0_f (new_AGEMA_signal_3211), .B1_t (new_AGEMA_signal_3212), .B1_f (new_AGEMA_signal_3213), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3635), .Z1_t (new_AGEMA_signal_3636), .Z1_f (new_AGEMA_signal_3637) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3635), .B1_t (new_AGEMA_signal_3636), .B1_f (new_AGEMA_signal_3637), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4057), .Z1_t (new_AGEMA_signal_4058), .Z1_f (new_AGEMA_signal_4059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4057), .A1_t (new_AGEMA_signal_4058), .A1_f (new_AGEMA_signal_4059), .B0_t (data_out_s0_t[6]), .B0_f (data_out_s0_f[6]), .B1_t (data_out_s1_t[6]), .B1_f (data_out_s1_f[6]), .Z0_t (data_out_s0_t[10]), .Z0_f (data_out_s0_f[10]), .Z1_t (data_out_s1_t[10]), .Z1_f (data_out_s1_f[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[7]), .A0_f (data_out_s0_f[7]), .A1_t (data_out_s1_t[7]), .A1_f (data_out_s1_f[7]), .B0_t (stateFF_inputPar[11]), .B0_f (new_AGEMA_signal_3214), .B1_t (new_AGEMA_signal_3215), .B1_f (new_AGEMA_signal_3216), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3638), .Z1_t (new_AGEMA_signal_3639), .Z1_f (new_AGEMA_signal_3640) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3638), .B1_t (new_AGEMA_signal_3639), .B1_f (new_AGEMA_signal_3640), .Z0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4060), .Z1_t (new_AGEMA_signal_4061), .Z1_f (new_AGEMA_signal_4062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4060), .A1_t (new_AGEMA_signal_4061), .A1_f (new_AGEMA_signal_4062), .B0_t (data_out_s0_t[7]), .B0_f (data_out_s0_f[7]), .B1_t (data_out_s1_t[7]), .B1_f (data_out_s1_f[7]), .Z0_t (data_out_s0_t[11]), .Z0_f (data_out_s0_f[11]), .Z1_t (data_out_s1_t[11]), .Z1_f (data_out_s1_f[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[8]), .A0_f (data_out_s0_f[8]), .A1_t (data_out_s1_t[8]), .A1_f (data_out_s1_f[8]), .B0_t (stateFF_inputPar[12]), .B0_f (new_AGEMA_signal_3217), .B1_t (new_AGEMA_signal_3218), .B1_f (new_AGEMA_signal_3219), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3641), .Z1_t (new_AGEMA_signal_3642), .Z1_f (new_AGEMA_signal_3643) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3641), .B1_t (new_AGEMA_signal_3642), .B1_f (new_AGEMA_signal_3643), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4063), .Z1_t (new_AGEMA_signal_4064), .Z1_f (new_AGEMA_signal_4065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4063), .A1_t (new_AGEMA_signal_4064), .A1_f (new_AGEMA_signal_4065), .B0_t (data_out_s0_t[8]), .B0_f (data_out_s0_f[8]), .B1_t (data_out_s1_t[8]), .B1_f (data_out_s1_f[8]), .Z0_t (data_out_s0_t[12]), .Z0_f (data_out_s0_f[12]), .Z1_t (data_out_s1_t[12]), .Z1_f (data_out_s1_f[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[9]), .A0_f (data_out_s0_f[9]), .A1_t (data_out_s1_t[9]), .A1_f (data_out_s1_f[9]), .B0_t (stateFF_inputPar[13]), .B0_f (new_AGEMA_signal_3220), .B1_t (new_AGEMA_signal_3221), .B1_f (new_AGEMA_signal_3222), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3644), .Z1_t (new_AGEMA_signal_3645), .Z1_f (new_AGEMA_signal_3646) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3644), .B1_t (new_AGEMA_signal_3645), .B1_f (new_AGEMA_signal_3646), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4066), .Z1_t (new_AGEMA_signal_4067), .Z1_f (new_AGEMA_signal_4068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4066), .A1_t (new_AGEMA_signal_4067), .A1_f (new_AGEMA_signal_4068), .B0_t (data_out_s0_t[9]), .B0_f (data_out_s0_f[9]), .B1_t (data_out_s1_t[9]), .B1_f (data_out_s1_f[9]), .Z0_t (data_out_s0_t[13]), .Z0_f (data_out_s0_f[13]), .Z1_t (data_out_s1_t[13]), .Z1_f (data_out_s1_f[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[10]), .A0_f (data_out_s0_f[10]), .A1_t (data_out_s1_t[10]), .A1_f (data_out_s1_f[10]), .B0_t (stateFF_inputPar[14]), .B0_f (new_AGEMA_signal_3223), .B1_t (new_AGEMA_signal_3224), .B1_f (new_AGEMA_signal_3225), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3647), .Z1_t (new_AGEMA_signal_3648), .Z1_f (new_AGEMA_signal_3649) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3647), .B1_t (new_AGEMA_signal_3648), .B1_f (new_AGEMA_signal_3649), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4069), .Z1_t (new_AGEMA_signal_4070), .Z1_f (new_AGEMA_signal_4071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4069), .A1_t (new_AGEMA_signal_4070), .A1_f (new_AGEMA_signal_4071), .B0_t (data_out_s0_t[10]), .B0_f (data_out_s0_f[10]), .B1_t (data_out_s1_t[10]), .B1_f (data_out_s1_f[10]), .Z0_t (data_out_s0_t[14]), .Z0_f (data_out_s0_f[14]), .Z1_t (data_out_s1_t[14]), .Z1_f (data_out_s1_f[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[11]), .A0_f (data_out_s0_f[11]), .A1_t (data_out_s1_t[11]), .A1_f (data_out_s1_f[11]), .B0_t (stateFF_inputPar[15]), .B0_f (new_AGEMA_signal_3226), .B1_t (new_AGEMA_signal_3227), .B1_f (new_AGEMA_signal_3228), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3650), .Z1_t (new_AGEMA_signal_3651), .Z1_f (new_AGEMA_signal_3652) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3650), .B1_t (new_AGEMA_signal_3651), .B1_f (new_AGEMA_signal_3652), .Z0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4072), .Z1_t (new_AGEMA_signal_4073), .Z1_f (new_AGEMA_signal_4074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4072), .A1_t (new_AGEMA_signal_4073), .A1_f (new_AGEMA_signal_4074), .B0_t (data_out_s0_t[11]), .B0_f (data_out_s0_f[11]), .B1_t (data_out_s1_t[11]), .B1_f (data_out_s1_f[11]), .Z0_t (data_out_s0_t[15]), .Z0_f (data_out_s0_f[15]), .Z1_t (data_out_s1_t[15]), .Z1_f (data_out_s1_f[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[12]), .A0_f (data_out_s0_f[12]), .A1_t (data_out_s1_t[12]), .A1_f (data_out_s1_f[12]), .B0_t (stateFF_inputPar[16]), .B0_f (new_AGEMA_signal_3229), .B1_t (new_AGEMA_signal_3230), .B1_f (new_AGEMA_signal_3231), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3653), .Z1_t (new_AGEMA_signal_3654), .Z1_f (new_AGEMA_signal_3655) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3653), .B1_t (new_AGEMA_signal_3654), .B1_f (new_AGEMA_signal_3655), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4075), .Z1_t (new_AGEMA_signal_4076), .Z1_f (new_AGEMA_signal_4077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4075), .A1_t (new_AGEMA_signal_4076), .A1_f (new_AGEMA_signal_4077), .B0_t (data_out_s0_t[12]), .B0_f (data_out_s0_f[12]), .B1_t (data_out_s1_t[12]), .B1_f (data_out_s1_f[12]), .Z0_t (data_out_s0_t[16]), .Z0_f (data_out_s0_f[16]), .Z1_t (data_out_s1_t[16]), .Z1_f (data_out_s1_f[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[13]), .A0_f (data_out_s0_f[13]), .A1_t (data_out_s1_t[13]), .A1_f (data_out_s1_f[13]), .B0_t (stateFF_inputPar[17]), .B0_f (new_AGEMA_signal_3232), .B1_t (new_AGEMA_signal_3233), .B1_f (new_AGEMA_signal_3234), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3656), .Z1_t (new_AGEMA_signal_3657), .Z1_f (new_AGEMA_signal_3658) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3656), .B1_t (new_AGEMA_signal_3657), .B1_f (new_AGEMA_signal_3658), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4078), .Z1_t (new_AGEMA_signal_4079), .Z1_f (new_AGEMA_signal_4080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4078), .A1_t (new_AGEMA_signal_4079), .A1_f (new_AGEMA_signal_4080), .B0_t (data_out_s0_t[13]), .B0_f (data_out_s0_f[13]), .B1_t (data_out_s1_t[13]), .B1_f (data_out_s1_f[13]), .Z0_t (data_out_s0_t[17]), .Z0_f (data_out_s0_f[17]), .Z1_t (data_out_s1_t[17]), .Z1_f (data_out_s1_f[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[14]), .A0_f (data_out_s0_f[14]), .A1_t (data_out_s1_t[14]), .A1_f (data_out_s1_f[14]), .B0_t (stateFF_inputPar[18]), .B0_f (new_AGEMA_signal_3235), .B1_t (new_AGEMA_signal_3236), .B1_f (new_AGEMA_signal_3237), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3659), .Z1_t (new_AGEMA_signal_3660), .Z1_f (new_AGEMA_signal_3661) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3659), .B1_t (new_AGEMA_signal_3660), .B1_f (new_AGEMA_signal_3661), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4081), .Z1_t (new_AGEMA_signal_4082), .Z1_f (new_AGEMA_signal_4083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4081), .A1_t (new_AGEMA_signal_4082), .A1_f (new_AGEMA_signal_4083), .B0_t (data_out_s0_t[14]), .B0_f (data_out_s0_f[14]), .B1_t (data_out_s1_t[14]), .B1_f (data_out_s1_f[14]), .Z0_t (data_out_s0_t[18]), .Z0_f (data_out_s0_f[18]), .Z1_t (data_out_s1_t[18]), .Z1_f (data_out_s1_f[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[15]), .A0_f (data_out_s0_f[15]), .A1_t (data_out_s1_t[15]), .A1_f (data_out_s1_f[15]), .B0_t (stateFF_inputPar[19]), .B0_f (new_AGEMA_signal_3238), .B1_t (new_AGEMA_signal_3239), .B1_f (new_AGEMA_signal_3240), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3662), .Z1_t (new_AGEMA_signal_3663), .Z1_f (new_AGEMA_signal_3664) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3662), .B1_t (new_AGEMA_signal_3663), .B1_f (new_AGEMA_signal_3664), .Z0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4084), .Z1_t (new_AGEMA_signal_4085), .Z1_f (new_AGEMA_signal_4086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4084), .A1_t (new_AGEMA_signal_4085), .A1_f (new_AGEMA_signal_4086), .B0_t (data_out_s0_t[15]), .B0_f (data_out_s0_f[15]), .B1_t (data_out_s1_t[15]), .B1_f (data_out_s1_f[15]), .Z0_t (data_out_s0_t[19]), .Z0_f (data_out_s0_f[19]), .Z1_t (data_out_s1_t[19]), .Z1_f (data_out_s1_f[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[16]), .A0_f (data_out_s0_f[16]), .A1_t (data_out_s1_t[16]), .A1_f (data_out_s1_f[16]), .B0_t (stateFF_inputPar[20]), .B0_f (new_AGEMA_signal_3241), .B1_t (new_AGEMA_signal_3242), .B1_f (new_AGEMA_signal_3243), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3665), .Z1_t (new_AGEMA_signal_3666), .Z1_f (new_AGEMA_signal_3667) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3665), .B1_t (new_AGEMA_signal_3666), .B1_f (new_AGEMA_signal_3667), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4087), .Z1_t (new_AGEMA_signal_4088), .Z1_f (new_AGEMA_signal_4089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4087), .A1_t (new_AGEMA_signal_4088), .A1_f (new_AGEMA_signal_4089), .B0_t (data_out_s0_t[16]), .B0_f (data_out_s0_f[16]), .B1_t (data_out_s1_t[16]), .B1_f (data_out_s1_f[16]), .Z0_t (data_out_s0_t[20]), .Z0_f (data_out_s0_f[20]), .Z1_t (data_out_s1_t[20]), .Z1_f (data_out_s1_f[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[17]), .A0_f (data_out_s0_f[17]), .A1_t (data_out_s1_t[17]), .A1_f (data_out_s1_f[17]), .B0_t (stateFF_inputPar[21]), .B0_f (new_AGEMA_signal_3244), .B1_t (new_AGEMA_signal_3245), .B1_f (new_AGEMA_signal_3246), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3668), .Z1_t (new_AGEMA_signal_3669), .Z1_f (new_AGEMA_signal_3670) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3668), .B1_t (new_AGEMA_signal_3669), .B1_f (new_AGEMA_signal_3670), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4090), .Z1_t (new_AGEMA_signal_4091), .Z1_f (new_AGEMA_signal_4092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4090), .A1_t (new_AGEMA_signal_4091), .A1_f (new_AGEMA_signal_4092), .B0_t (data_out_s0_t[17]), .B0_f (data_out_s0_f[17]), .B1_t (data_out_s1_t[17]), .B1_f (data_out_s1_f[17]), .Z0_t (data_out_s0_t[21]), .Z0_f (data_out_s0_f[21]), .Z1_t (data_out_s1_t[21]), .Z1_f (data_out_s1_f[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[18]), .A0_f (data_out_s0_f[18]), .A1_t (data_out_s1_t[18]), .A1_f (data_out_s1_f[18]), .B0_t (stateFF_inputPar[22]), .B0_f (new_AGEMA_signal_3247), .B1_t (new_AGEMA_signal_3248), .B1_f (new_AGEMA_signal_3249), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3671), .Z1_t (new_AGEMA_signal_3672), .Z1_f (new_AGEMA_signal_3673) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3671), .B1_t (new_AGEMA_signal_3672), .B1_f (new_AGEMA_signal_3673), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4093), .Z1_t (new_AGEMA_signal_4094), .Z1_f (new_AGEMA_signal_4095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4093), .A1_t (new_AGEMA_signal_4094), .A1_f (new_AGEMA_signal_4095), .B0_t (data_out_s0_t[18]), .B0_f (data_out_s0_f[18]), .B1_t (data_out_s1_t[18]), .B1_f (data_out_s1_f[18]), .Z0_t (data_out_s0_t[22]), .Z0_f (data_out_s0_f[22]), .Z1_t (data_out_s1_t[22]), .Z1_f (data_out_s1_f[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[19]), .A0_f (data_out_s0_f[19]), .A1_t (data_out_s1_t[19]), .A1_f (data_out_s1_f[19]), .B0_t (stateFF_inputPar[23]), .B0_f (new_AGEMA_signal_3250), .B1_t (new_AGEMA_signal_3251), .B1_f (new_AGEMA_signal_3252), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3674), .Z1_t (new_AGEMA_signal_3675), .Z1_f (new_AGEMA_signal_3676) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3674), .B1_t (new_AGEMA_signal_3675), .B1_f (new_AGEMA_signal_3676), .Z0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4096), .Z1_t (new_AGEMA_signal_4097), .Z1_f (new_AGEMA_signal_4098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4096), .A1_t (new_AGEMA_signal_4097), .A1_f (new_AGEMA_signal_4098), .B0_t (data_out_s0_t[19]), .B0_f (data_out_s0_f[19]), .B1_t (data_out_s1_t[19]), .B1_f (data_out_s1_f[19]), .Z0_t (data_out_s0_t[23]), .Z0_f (data_out_s0_f[23]), .Z1_t (data_out_s1_t[23]), .Z1_f (data_out_s1_f[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[20]), .A0_f (data_out_s0_f[20]), .A1_t (data_out_s1_t[20]), .A1_f (data_out_s1_f[20]), .B0_t (stateFF_inputPar[24]), .B0_f (new_AGEMA_signal_3253), .B1_t (new_AGEMA_signal_3254), .B1_f (new_AGEMA_signal_3255), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3677), .Z1_t (new_AGEMA_signal_3678), .Z1_f (new_AGEMA_signal_3679) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3677), .B1_t (new_AGEMA_signal_3678), .B1_f (new_AGEMA_signal_3679), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4099), .Z1_t (new_AGEMA_signal_4100), .Z1_f (new_AGEMA_signal_4101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4099), .A1_t (new_AGEMA_signal_4100), .A1_f (new_AGEMA_signal_4101), .B0_t (data_out_s0_t[20]), .B0_f (data_out_s0_f[20]), .B1_t (data_out_s1_t[20]), .B1_f (data_out_s1_f[20]), .Z0_t (data_out_s0_t[24]), .Z0_f (data_out_s0_f[24]), .Z1_t (data_out_s1_t[24]), .Z1_f (data_out_s1_f[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[21]), .A0_f (data_out_s0_f[21]), .A1_t (data_out_s1_t[21]), .A1_f (data_out_s1_f[21]), .B0_t (stateFF_inputPar[25]), .B0_f (new_AGEMA_signal_3256), .B1_t (new_AGEMA_signal_3257), .B1_f (new_AGEMA_signal_3258), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3680), .Z1_t (new_AGEMA_signal_3681), .Z1_f (new_AGEMA_signal_3682) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3680), .B1_t (new_AGEMA_signal_3681), .B1_f (new_AGEMA_signal_3682), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4102), .Z1_t (new_AGEMA_signal_4103), .Z1_f (new_AGEMA_signal_4104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4102), .A1_t (new_AGEMA_signal_4103), .A1_f (new_AGEMA_signal_4104), .B0_t (data_out_s0_t[21]), .B0_f (data_out_s0_f[21]), .B1_t (data_out_s1_t[21]), .B1_f (data_out_s1_f[21]), .Z0_t (data_out_s0_t[25]), .Z0_f (data_out_s0_f[25]), .Z1_t (data_out_s1_t[25]), .Z1_f (data_out_s1_f[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[22]), .A0_f (data_out_s0_f[22]), .A1_t (data_out_s1_t[22]), .A1_f (data_out_s1_f[22]), .B0_t (stateFF_inputPar[26]), .B0_f (new_AGEMA_signal_3259), .B1_t (new_AGEMA_signal_3260), .B1_f (new_AGEMA_signal_3261), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3683), .Z1_t (new_AGEMA_signal_3684), .Z1_f (new_AGEMA_signal_3685) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3683), .B1_t (new_AGEMA_signal_3684), .B1_f (new_AGEMA_signal_3685), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4105), .Z1_t (new_AGEMA_signal_4106), .Z1_f (new_AGEMA_signal_4107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4105), .A1_t (new_AGEMA_signal_4106), .A1_f (new_AGEMA_signal_4107), .B0_t (data_out_s0_t[22]), .B0_f (data_out_s0_f[22]), .B1_t (data_out_s1_t[22]), .B1_f (data_out_s1_f[22]), .Z0_t (data_out_s0_t[26]), .Z0_f (data_out_s0_f[26]), .Z1_t (data_out_s1_t[26]), .Z1_f (data_out_s1_f[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[23]), .A0_f (data_out_s0_f[23]), .A1_t (data_out_s1_t[23]), .A1_f (data_out_s1_f[23]), .B0_t (stateFF_inputPar[27]), .B0_f (new_AGEMA_signal_3262), .B1_t (new_AGEMA_signal_3263), .B1_f (new_AGEMA_signal_3264), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3686), .Z1_t (new_AGEMA_signal_3687), .Z1_f (new_AGEMA_signal_3688) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3686), .B1_t (new_AGEMA_signal_3687), .B1_f (new_AGEMA_signal_3688), .Z0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4108), .Z1_t (new_AGEMA_signal_4109), .Z1_f (new_AGEMA_signal_4110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4108), .A1_t (new_AGEMA_signal_4109), .A1_f (new_AGEMA_signal_4110), .B0_t (data_out_s0_t[23]), .B0_f (data_out_s0_f[23]), .B1_t (data_out_s1_t[23]), .B1_f (data_out_s1_f[23]), .Z0_t (data_out_s0_t[27]), .Z0_f (data_out_s0_f[27]), .Z1_t (data_out_s1_t[27]), .Z1_f (data_out_s1_f[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[24]), .A0_f (data_out_s0_f[24]), .A1_t (data_out_s1_t[24]), .A1_f (data_out_s1_f[24]), .B0_t (stateFF_inputPar[28]), .B0_f (new_AGEMA_signal_3265), .B1_t (new_AGEMA_signal_3266), .B1_f (new_AGEMA_signal_3267), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3689), .Z1_t (new_AGEMA_signal_3690), .Z1_f (new_AGEMA_signal_3691) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3689), .B1_t (new_AGEMA_signal_3690), .B1_f (new_AGEMA_signal_3691), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4111), .Z1_t (new_AGEMA_signal_4112), .Z1_f (new_AGEMA_signal_4113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4111), .A1_t (new_AGEMA_signal_4112), .A1_f (new_AGEMA_signal_4113), .B0_t (data_out_s0_t[24]), .B0_f (data_out_s0_f[24]), .B1_t (data_out_s1_t[24]), .B1_f (data_out_s1_f[24]), .Z0_t (data_out_s0_t[28]), .Z0_f (data_out_s0_f[28]), .Z1_t (data_out_s1_t[28]), .Z1_f (data_out_s1_f[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[25]), .A0_f (data_out_s0_f[25]), .A1_t (data_out_s1_t[25]), .A1_f (data_out_s1_f[25]), .B0_t (stateFF_inputPar[29]), .B0_f (new_AGEMA_signal_3268), .B1_t (new_AGEMA_signal_3269), .B1_f (new_AGEMA_signal_3270), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3692), .Z1_t (new_AGEMA_signal_3693), .Z1_f (new_AGEMA_signal_3694) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3692), .B1_t (new_AGEMA_signal_3693), .B1_f (new_AGEMA_signal_3694), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4114), .Z1_t (new_AGEMA_signal_4115), .Z1_f (new_AGEMA_signal_4116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4114), .A1_t (new_AGEMA_signal_4115), .A1_f (new_AGEMA_signal_4116), .B0_t (data_out_s0_t[25]), .B0_f (data_out_s0_f[25]), .B1_t (data_out_s1_t[25]), .B1_f (data_out_s1_f[25]), .Z0_t (data_out_s0_t[29]), .Z0_f (data_out_s0_f[29]), .Z1_t (data_out_s1_t[29]), .Z1_f (data_out_s1_f[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[26]), .A0_f (data_out_s0_f[26]), .A1_t (data_out_s1_t[26]), .A1_f (data_out_s1_f[26]), .B0_t (stateFF_inputPar[30]), .B0_f (new_AGEMA_signal_3271), .B1_t (new_AGEMA_signal_3272), .B1_f (new_AGEMA_signal_3273), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3695), .Z1_t (new_AGEMA_signal_3696), .Z1_f (new_AGEMA_signal_3697) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3695), .B1_t (new_AGEMA_signal_3696), .B1_f (new_AGEMA_signal_3697), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4117), .Z1_t (new_AGEMA_signal_4118), .Z1_f (new_AGEMA_signal_4119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4117), .A1_t (new_AGEMA_signal_4118), .A1_f (new_AGEMA_signal_4119), .B0_t (data_out_s0_t[26]), .B0_f (data_out_s0_f[26]), .B1_t (data_out_s1_t[26]), .B1_f (data_out_s1_f[26]), .Z0_t (data_out_s0_t[30]), .Z0_f (data_out_s0_f[30]), .Z1_t (data_out_s1_t[30]), .Z1_f (data_out_s1_f[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[27]), .A0_f (data_out_s0_f[27]), .A1_t (data_out_s1_t[27]), .A1_f (data_out_s1_f[27]), .B0_t (stateFF_inputPar[31]), .B0_f (new_AGEMA_signal_3274), .B1_t (new_AGEMA_signal_3275), .B1_f (new_AGEMA_signal_3276), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3698), .Z1_t (new_AGEMA_signal_3699), .Z1_f (new_AGEMA_signal_3700) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3698), .B1_t (new_AGEMA_signal_3699), .B1_f (new_AGEMA_signal_3700), .Z0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4120), .Z1_t (new_AGEMA_signal_4121), .Z1_f (new_AGEMA_signal_4122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4120), .A1_t (new_AGEMA_signal_4121), .A1_f (new_AGEMA_signal_4122), .B0_t (data_out_s0_t[27]), .B0_f (data_out_s0_f[27]), .B1_t (data_out_s1_t[27]), .B1_f (data_out_s1_f[27]), .Z0_t (data_out_s0_t[31]), .Z0_f (data_out_s0_f[31]), .Z1_t (data_out_s1_t[31]), .Z1_f (data_out_s1_f[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[28]), .A0_f (data_out_s0_f[28]), .A1_t (data_out_s1_t[28]), .A1_f (data_out_s1_f[28]), .B0_t (stateFF_inputPar[32]), .B0_f (new_AGEMA_signal_3277), .B1_t (new_AGEMA_signal_3278), .B1_f (new_AGEMA_signal_3279), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3701), .Z1_t (new_AGEMA_signal_3702), .Z1_f (new_AGEMA_signal_3703) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3701), .B1_t (new_AGEMA_signal_3702), .B1_f (new_AGEMA_signal_3703), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4123), .Z1_t (new_AGEMA_signal_4124), .Z1_f (new_AGEMA_signal_4125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4123), .A1_t (new_AGEMA_signal_4124), .A1_f (new_AGEMA_signal_4125), .B0_t (data_out_s0_t[28]), .B0_f (data_out_s0_f[28]), .B1_t (data_out_s1_t[28]), .B1_f (data_out_s1_f[28]), .Z0_t (data_out_s0_t[32]), .Z0_f (data_out_s0_f[32]), .Z1_t (data_out_s1_t[32]), .Z1_f (data_out_s1_f[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[29]), .A0_f (data_out_s0_f[29]), .A1_t (data_out_s1_t[29]), .A1_f (data_out_s1_f[29]), .B0_t (stateFF_inputPar[33]), .B0_f (new_AGEMA_signal_3280), .B1_t (new_AGEMA_signal_3281), .B1_f (new_AGEMA_signal_3282), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3704), .Z1_t (new_AGEMA_signal_3705), .Z1_f (new_AGEMA_signal_3706) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3704), .B1_t (new_AGEMA_signal_3705), .B1_f (new_AGEMA_signal_3706), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4126), .Z1_t (new_AGEMA_signal_4127), .Z1_f (new_AGEMA_signal_4128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4126), .A1_t (new_AGEMA_signal_4127), .A1_f (new_AGEMA_signal_4128), .B0_t (data_out_s0_t[29]), .B0_f (data_out_s0_f[29]), .B1_t (data_out_s1_t[29]), .B1_f (data_out_s1_f[29]), .Z0_t (data_out_s0_t[33]), .Z0_f (data_out_s0_f[33]), .Z1_t (data_out_s1_t[33]), .Z1_f (data_out_s1_f[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[30]), .A0_f (data_out_s0_f[30]), .A1_t (data_out_s1_t[30]), .A1_f (data_out_s1_f[30]), .B0_t (stateFF_inputPar[34]), .B0_f (new_AGEMA_signal_3283), .B1_t (new_AGEMA_signal_3284), .B1_f (new_AGEMA_signal_3285), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3707), .Z1_t (new_AGEMA_signal_3708), .Z1_f (new_AGEMA_signal_3709) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3707), .B1_t (new_AGEMA_signal_3708), .B1_f (new_AGEMA_signal_3709), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4129), .Z1_t (new_AGEMA_signal_4130), .Z1_f (new_AGEMA_signal_4131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4129), .A1_t (new_AGEMA_signal_4130), .A1_f (new_AGEMA_signal_4131), .B0_t (data_out_s0_t[30]), .B0_f (data_out_s0_f[30]), .B1_t (data_out_s1_t[30]), .B1_f (data_out_s1_f[30]), .Z0_t (data_out_s0_t[34]), .Z0_f (data_out_s0_f[34]), .Z1_t (data_out_s1_t[34]), .Z1_f (data_out_s1_f[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[31]), .A0_f (data_out_s0_f[31]), .A1_t (data_out_s1_t[31]), .A1_f (data_out_s1_f[31]), .B0_t (stateFF_inputPar[35]), .B0_f (new_AGEMA_signal_3286), .B1_t (new_AGEMA_signal_3287), .B1_f (new_AGEMA_signal_3288), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3710), .Z1_t (new_AGEMA_signal_3711), .Z1_f (new_AGEMA_signal_3712) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3710), .B1_t (new_AGEMA_signal_3711), .B1_f (new_AGEMA_signal_3712), .Z0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4132), .Z1_t (new_AGEMA_signal_4133), .Z1_f (new_AGEMA_signal_4134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4132), .A1_t (new_AGEMA_signal_4133), .A1_f (new_AGEMA_signal_4134), .B0_t (data_out_s0_t[31]), .B0_f (data_out_s0_f[31]), .B1_t (data_out_s1_t[31]), .B1_f (data_out_s1_f[31]), .Z0_t (data_out_s0_t[35]), .Z0_f (data_out_s0_f[35]), .Z1_t (data_out_s1_t[35]), .Z1_f (data_out_s1_f[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[32]), .A0_f (data_out_s0_f[32]), .A1_t (data_out_s1_t[32]), .A1_f (data_out_s1_f[32]), .B0_t (stateFF_inputPar[36]), .B0_f (new_AGEMA_signal_3289), .B1_t (new_AGEMA_signal_3290), .B1_f (new_AGEMA_signal_3291), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3713), .Z1_t (new_AGEMA_signal_3714), .Z1_f (new_AGEMA_signal_3715) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3713), .B1_t (new_AGEMA_signal_3714), .B1_f (new_AGEMA_signal_3715), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4135), .Z1_t (new_AGEMA_signal_4136), .Z1_f (new_AGEMA_signal_4137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4135), .A1_t (new_AGEMA_signal_4136), .A1_f (new_AGEMA_signal_4137), .B0_t (data_out_s0_t[32]), .B0_f (data_out_s0_f[32]), .B1_t (data_out_s1_t[32]), .B1_f (data_out_s1_f[32]), .Z0_t (data_out_s0_t[36]), .Z0_f (data_out_s0_f[36]), .Z1_t (data_out_s1_t[36]), .Z1_f (data_out_s1_f[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[33]), .A0_f (data_out_s0_f[33]), .A1_t (data_out_s1_t[33]), .A1_f (data_out_s1_f[33]), .B0_t (stateFF_inputPar[37]), .B0_f (new_AGEMA_signal_3292), .B1_t (new_AGEMA_signal_3293), .B1_f (new_AGEMA_signal_3294), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3716), .Z1_t (new_AGEMA_signal_3717), .Z1_f (new_AGEMA_signal_3718) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3716), .B1_t (new_AGEMA_signal_3717), .B1_f (new_AGEMA_signal_3718), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4138), .Z1_t (new_AGEMA_signal_4139), .Z1_f (new_AGEMA_signal_4140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4138), .A1_t (new_AGEMA_signal_4139), .A1_f (new_AGEMA_signal_4140), .B0_t (data_out_s0_t[33]), .B0_f (data_out_s0_f[33]), .B1_t (data_out_s1_t[33]), .B1_f (data_out_s1_f[33]), .Z0_t (data_out_s0_t[37]), .Z0_f (data_out_s0_f[37]), .Z1_t (data_out_s1_t[37]), .Z1_f (data_out_s1_f[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[34]), .A0_f (data_out_s0_f[34]), .A1_t (data_out_s1_t[34]), .A1_f (data_out_s1_f[34]), .B0_t (stateFF_inputPar[38]), .B0_f (new_AGEMA_signal_3295), .B1_t (new_AGEMA_signal_3296), .B1_f (new_AGEMA_signal_3297), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3719), .Z1_t (new_AGEMA_signal_3720), .Z1_f (new_AGEMA_signal_3721) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3719), .B1_t (new_AGEMA_signal_3720), .B1_f (new_AGEMA_signal_3721), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4141), .Z1_t (new_AGEMA_signal_4142), .Z1_f (new_AGEMA_signal_4143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4141), .A1_t (new_AGEMA_signal_4142), .A1_f (new_AGEMA_signal_4143), .B0_t (data_out_s0_t[34]), .B0_f (data_out_s0_f[34]), .B1_t (data_out_s1_t[34]), .B1_f (data_out_s1_f[34]), .Z0_t (data_out_s0_t[38]), .Z0_f (data_out_s0_f[38]), .Z1_t (data_out_s1_t[38]), .Z1_f (data_out_s1_f[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[35]), .A0_f (data_out_s0_f[35]), .A1_t (data_out_s1_t[35]), .A1_f (data_out_s1_f[35]), .B0_t (stateFF_inputPar[39]), .B0_f (new_AGEMA_signal_3298), .B1_t (new_AGEMA_signal_3299), .B1_f (new_AGEMA_signal_3300), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3722), .Z1_t (new_AGEMA_signal_3723), .Z1_f (new_AGEMA_signal_3724) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3722), .B1_t (new_AGEMA_signal_3723), .B1_f (new_AGEMA_signal_3724), .Z0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4144), .Z1_t (new_AGEMA_signal_4145), .Z1_f (new_AGEMA_signal_4146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4144), .A1_t (new_AGEMA_signal_4145), .A1_f (new_AGEMA_signal_4146), .B0_t (data_out_s0_t[35]), .B0_f (data_out_s0_f[35]), .B1_t (data_out_s1_t[35]), .B1_f (data_out_s1_f[35]), .Z0_t (data_out_s0_t[39]), .Z0_f (data_out_s0_f[39]), .Z1_t (data_out_s1_t[39]), .Z1_f (data_out_s1_f[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[36]), .A0_f (data_out_s0_f[36]), .A1_t (data_out_s1_t[36]), .A1_f (data_out_s1_f[36]), .B0_t (stateFF_inputPar[40]), .B0_f (new_AGEMA_signal_3301), .B1_t (new_AGEMA_signal_3302), .B1_f (new_AGEMA_signal_3303), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3725), .Z1_t (new_AGEMA_signal_3726), .Z1_f (new_AGEMA_signal_3727) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3725), .B1_t (new_AGEMA_signal_3726), .B1_f (new_AGEMA_signal_3727), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4147), .Z1_t (new_AGEMA_signal_4148), .Z1_f (new_AGEMA_signal_4149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4147), .A1_t (new_AGEMA_signal_4148), .A1_f (new_AGEMA_signal_4149), .B0_t (data_out_s0_t[36]), .B0_f (data_out_s0_f[36]), .B1_t (data_out_s1_t[36]), .B1_f (data_out_s1_f[36]), .Z0_t (data_out_s0_t[40]), .Z0_f (data_out_s0_f[40]), .Z1_t (data_out_s1_t[40]), .Z1_f (data_out_s1_f[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[37]), .A0_f (data_out_s0_f[37]), .A1_t (data_out_s1_t[37]), .A1_f (data_out_s1_f[37]), .B0_t (stateFF_inputPar[41]), .B0_f (new_AGEMA_signal_3304), .B1_t (new_AGEMA_signal_3305), .B1_f (new_AGEMA_signal_3306), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3728), .Z1_t (new_AGEMA_signal_3729), .Z1_f (new_AGEMA_signal_3730) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3728), .B1_t (new_AGEMA_signal_3729), .B1_f (new_AGEMA_signal_3730), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4150), .Z1_t (new_AGEMA_signal_4151), .Z1_f (new_AGEMA_signal_4152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4150), .A1_t (new_AGEMA_signal_4151), .A1_f (new_AGEMA_signal_4152), .B0_t (data_out_s0_t[37]), .B0_f (data_out_s0_f[37]), .B1_t (data_out_s1_t[37]), .B1_f (data_out_s1_f[37]), .Z0_t (data_out_s0_t[41]), .Z0_f (data_out_s0_f[41]), .Z1_t (data_out_s1_t[41]), .Z1_f (data_out_s1_f[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[38]), .A0_f (data_out_s0_f[38]), .A1_t (data_out_s1_t[38]), .A1_f (data_out_s1_f[38]), .B0_t (stateFF_inputPar[42]), .B0_f (new_AGEMA_signal_3307), .B1_t (new_AGEMA_signal_3308), .B1_f (new_AGEMA_signal_3309), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3731), .Z1_t (new_AGEMA_signal_3732), .Z1_f (new_AGEMA_signal_3733) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3731), .B1_t (new_AGEMA_signal_3732), .B1_f (new_AGEMA_signal_3733), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4153), .Z1_t (new_AGEMA_signal_4154), .Z1_f (new_AGEMA_signal_4155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4153), .A1_t (new_AGEMA_signal_4154), .A1_f (new_AGEMA_signal_4155), .B0_t (data_out_s0_t[38]), .B0_f (data_out_s0_f[38]), .B1_t (data_out_s1_t[38]), .B1_f (data_out_s1_f[38]), .Z0_t (data_out_s0_t[42]), .Z0_f (data_out_s0_f[42]), .Z1_t (data_out_s1_t[42]), .Z1_f (data_out_s1_f[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[39]), .A0_f (data_out_s0_f[39]), .A1_t (data_out_s1_t[39]), .A1_f (data_out_s1_f[39]), .B0_t (stateFF_inputPar[43]), .B0_f (new_AGEMA_signal_3310), .B1_t (new_AGEMA_signal_3311), .B1_f (new_AGEMA_signal_3312), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3734), .Z1_t (new_AGEMA_signal_3735), .Z1_f (new_AGEMA_signal_3736) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3734), .B1_t (new_AGEMA_signal_3735), .B1_f (new_AGEMA_signal_3736), .Z0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4156), .Z1_t (new_AGEMA_signal_4157), .Z1_f (new_AGEMA_signal_4158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4156), .A1_t (new_AGEMA_signal_4157), .A1_f (new_AGEMA_signal_4158), .B0_t (data_out_s0_t[39]), .B0_f (data_out_s0_f[39]), .B1_t (data_out_s1_t[39]), .B1_f (data_out_s1_f[39]), .Z0_t (data_out_s0_t[43]), .Z0_f (data_out_s0_f[43]), .Z1_t (data_out_s1_t[43]), .Z1_f (data_out_s1_f[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[40]), .A0_f (data_out_s0_f[40]), .A1_t (data_out_s1_t[40]), .A1_f (data_out_s1_f[40]), .B0_t (stateFF_inputPar[44]), .B0_f (new_AGEMA_signal_3313), .B1_t (new_AGEMA_signal_3314), .B1_f (new_AGEMA_signal_3315), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3737), .Z1_t (new_AGEMA_signal_3738), .Z1_f (new_AGEMA_signal_3739) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3737), .B1_t (new_AGEMA_signal_3738), .B1_f (new_AGEMA_signal_3739), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4159), .Z1_t (new_AGEMA_signal_4160), .Z1_f (new_AGEMA_signal_4161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4159), .A1_t (new_AGEMA_signal_4160), .A1_f (new_AGEMA_signal_4161), .B0_t (data_out_s0_t[40]), .B0_f (data_out_s0_f[40]), .B1_t (data_out_s1_t[40]), .B1_f (data_out_s1_f[40]), .Z0_t (data_out_s0_t[44]), .Z0_f (data_out_s0_f[44]), .Z1_t (data_out_s1_t[44]), .Z1_f (data_out_s1_f[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[41]), .A0_f (data_out_s0_f[41]), .A1_t (data_out_s1_t[41]), .A1_f (data_out_s1_f[41]), .B0_t (stateFF_inputPar[45]), .B0_f (new_AGEMA_signal_3316), .B1_t (new_AGEMA_signal_3317), .B1_f (new_AGEMA_signal_3318), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3740), .Z1_t (new_AGEMA_signal_3741), .Z1_f (new_AGEMA_signal_3742) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3740), .B1_t (new_AGEMA_signal_3741), .B1_f (new_AGEMA_signal_3742), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4162), .Z1_t (new_AGEMA_signal_4163), .Z1_f (new_AGEMA_signal_4164) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4162), .A1_t (new_AGEMA_signal_4163), .A1_f (new_AGEMA_signal_4164), .B0_t (data_out_s0_t[41]), .B0_f (data_out_s0_f[41]), .B1_t (data_out_s1_t[41]), .B1_f (data_out_s1_f[41]), .Z0_t (data_out_s0_t[45]), .Z0_f (data_out_s0_f[45]), .Z1_t (data_out_s1_t[45]), .Z1_f (data_out_s1_f[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[42]), .A0_f (data_out_s0_f[42]), .A1_t (data_out_s1_t[42]), .A1_f (data_out_s1_f[42]), .B0_t (stateFF_inputPar[46]), .B0_f (new_AGEMA_signal_3319), .B1_t (new_AGEMA_signal_3320), .B1_f (new_AGEMA_signal_3321), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3743), .Z1_t (new_AGEMA_signal_3744), .Z1_f (new_AGEMA_signal_3745) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3743), .B1_t (new_AGEMA_signal_3744), .B1_f (new_AGEMA_signal_3745), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4165), .Z1_t (new_AGEMA_signal_4166), .Z1_f (new_AGEMA_signal_4167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4165), .A1_t (new_AGEMA_signal_4166), .A1_f (new_AGEMA_signal_4167), .B0_t (data_out_s0_t[42]), .B0_f (data_out_s0_f[42]), .B1_t (data_out_s1_t[42]), .B1_f (data_out_s1_f[42]), .Z0_t (data_out_s0_t[46]), .Z0_f (data_out_s0_f[46]), .Z1_t (data_out_s1_t[46]), .Z1_f (data_out_s1_f[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[43]), .A0_f (data_out_s0_f[43]), .A1_t (data_out_s1_t[43]), .A1_f (data_out_s1_f[43]), .B0_t (stateFF_inputPar[47]), .B0_f (new_AGEMA_signal_3322), .B1_t (new_AGEMA_signal_3323), .B1_f (new_AGEMA_signal_3324), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3746), .Z1_t (new_AGEMA_signal_3747), .Z1_f (new_AGEMA_signal_3748) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3746), .B1_t (new_AGEMA_signal_3747), .B1_f (new_AGEMA_signal_3748), .Z0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4168), .Z1_t (new_AGEMA_signal_4169), .Z1_f (new_AGEMA_signal_4170) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4168), .A1_t (new_AGEMA_signal_4169), .A1_f (new_AGEMA_signal_4170), .B0_t (data_out_s0_t[43]), .B0_f (data_out_s0_f[43]), .B1_t (data_out_s1_t[43]), .B1_f (data_out_s1_f[43]), .Z0_t (data_out_s0_t[47]), .Z0_f (data_out_s0_f[47]), .Z1_t (data_out_s1_t[47]), .Z1_f (data_out_s1_f[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[44]), .A0_f (data_out_s0_f[44]), .A1_t (data_out_s1_t[44]), .A1_f (data_out_s1_f[44]), .B0_t (stateFF_inputPar[48]), .B0_f (new_AGEMA_signal_3325), .B1_t (new_AGEMA_signal_3326), .B1_f (new_AGEMA_signal_3327), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3749), .Z1_t (new_AGEMA_signal_3750), .Z1_f (new_AGEMA_signal_3751) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3749), .B1_t (new_AGEMA_signal_3750), .B1_f (new_AGEMA_signal_3751), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4171), .Z1_t (new_AGEMA_signal_4172), .Z1_f (new_AGEMA_signal_4173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4171), .A1_t (new_AGEMA_signal_4172), .A1_f (new_AGEMA_signal_4173), .B0_t (data_out_s0_t[44]), .B0_f (data_out_s0_f[44]), .B1_t (data_out_s1_t[44]), .B1_f (data_out_s1_f[44]), .Z0_t (data_out_s0_t[48]), .Z0_f (data_out_s0_f[48]), .Z1_t (data_out_s1_t[48]), .Z1_f (data_out_s1_f[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[45]), .A0_f (data_out_s0_f[45]), .A1_t (data_out_s1_t[45]), .A1_f (data_out_s1_f[45]), .B0_t (stateFF_inputPar[49]), .B0_f (new_AGEMA_signal_3328), .B1_t (new_AGEMA_signal_3329), .B1_f (new_AGEMA_signal_3330), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3752), .Z1_t (new_AGEMA_signal_3753), .Z1_f (new_AGEMA_signal_3754) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3752), .B1_t (new_AGEMA_signal_3753), .B1_f (new_AGEMA_signal_3754), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4174), .Z1_t (new_AGEMA_signal_4175), .Z1_f (new_AGEMA_signal_4176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4174), .A1_t (new_AGEMA_signal_4175), .A1_f (new_AGEMA_signal_4176), .B0_t (data_out_s0_t[45]), .B0_f (data_out_s0_f[45]), .B1_t (data_out_s1_t[45]), .B1_f (data_out_s1_f[45]), .Z0_t (data_out_s0_t[49]), .Z0_f (data_out_s0_f[49]), .Z1_t (data_out_s1_t[49]), .Z1_f (data_out_s1_f[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[46]), .A0_f (data_out_s0_f[46]), .A1_t (data_out_s1_t[46]), .A1_f (data_out_s1_f[46]), .B0_t (stateFF_inputPar[50]), .B0_f (new_AGEMA_signal_3331), .B1_t (new_AGEMA_signal_3332), .B1_f (new_AGEMA_signal_3333), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3755), .Z1_t (new_AGEMA_signal_3756), .Z1_f (new_AGEMA_signal_3757) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3755), .B1_t (new_AGEMA_signal_3756), .B1_f (new_AGEMA_signal_3757), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4177), .Z1_t (new_AGEMA_signal_4178), .Z1_f (new_AGEMA_signal_4179) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4177), .A1_t (new_AGEMA_signal_4178), .A1_f (new_AGEMA_signal_4179), .B0_t (data_out_s0_t[46]), .B0_f (data_out_s0_f[46]), .B1_t (data_out_s1_t[46]), .B1_f (data_out_s1_f[46]), .Z0_t (data_out_s0_t[50]), .Z0_f (data_out_s0_f[50]), .Z1_t (data_out_s1_t[50]), .Z1_f (data_out_s1_f[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[47]), .A0_f (data_out_s0_f[47]), .A1_t (data_out_s1_t[47]), .A1_f (data_out_s1_f[47]), .B0_t (stateFF_inputPar[51]), .B0_f (new_AGEMA_signal_3334), .B1_t (new_AGEMA_signal_3335), .B1_f (new_AGEMA_signal_3336), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3758), .Z1_t (new_AGEMA_signal_3759), .Z1_f (new_AGEMA_signal_3760) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3758), .B1_t (new_AGEMA_signal_3759), .B1_f (new_AGEMA_signal_3760), .Z0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4180), .Z1_t (new_AGEMA_signal_4181), .Z1_f (new_AGEMA_signal_4182) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4180), .A1_t (new_AGEMA_signal_4181), .A1_f (new_AGEMA_signal_4182), .B0_t (data_out_s0_t[47]), .B0_f (data_out_s0_f[47]), .B1_t (data_out_s1_t[47]), .B1_f (data_out_s1_f[47]), .Z0_t (data_out_s0_t[51]), .Z0_f (data_out_s0_f[51]), .Z1_t (data_out_s1_t[51]), .Z1_f (data_out_s1_f[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[48]), .A0_f (data_out_s0_f[48]), .A1_t (data_out_s1_t[48]), .A1_f (data_out_s1_f[48]), .B0_t (stateFF_inputPar[52]), .B0_f (new_AGEMA_signal_3337), .B1_t (new_AGEMA_signal_3338), .B1_f (new_AGEMA_signal_3339), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3761), .Z1_t (new_AGEMA_signal_3762), .Z1_f (new_AGEMA_signal_3763) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3761), .B1_t (new_AGEMA_signal_3762), .B1_f (new_AGEMA_signal_3763), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4183), .Z1_t (new_AGEMA_signal_4184), .Z1_f (new_AGEMA_signal_4185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4183), .A1_t (new_AGEMA_signal_4184), .A1_f (new_AGEMA_signal_4185), .B0_t (data_out_s0_t[48]), .B0_f (data_out_s0_f[48]), .B1_t (data_out_s1_t[48]), .B1_f (data_out_s1_f[48]), .Z0_t (data_out_s0_t[52]), .Z0_f (data_out_s0_f[52]), .Z1_t (data_out_s1_t[52]), .Z1_f (data_out_s1_f[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[49]), .A0_f (data_out_s0_f[49]), .A1_t (data_out_s1_t[49]), .A1_f (data_out_s1_f[49]), .B0_t (stateFF_inputPar[53]), .B0_f (new_AGEMA_signal_3340), .B1_t (new_AGEMA_signal_3341), .B1_f (new_AGEMA_signal_3342), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3764), .Z1_t (new_AGEMA_signal_3765), .Z1_f (new_AGEMA_signal_3766) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3764), .B1_t (new_AGEMA_signal_3765), .B1_f (new_AGEMA_signal_3766), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4186), .Z1_t (new_AGEMA_signal_4187), .Z1_f (new_AGEMA_signal_4188) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4186), .A1_t (new_AGEMA_signal_4187), .A1_f (new_AGEMA_signal_4188), .B0_t (data_out_s0_t[49]), .B0_f (data_out_s0_f[49]), .B1_t (data_out_s1_t[49]), .B1_f (data_out_s1_f[49]), .Z0_t (data_out_s0_t[53]), .Z0_f (data_out_s0_f[53]), .Z1_t (data_out_s1_t[53]), .Z1_f (data_out_s1_f[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[50]), .A0_f (data_out_s0_f[50]), .A1_t (data_out_s1_t[50]), .A1_f (data_out_s1_f[50]), .B0_t (stateFF_inputPar[54]), .B0_f (new_AGEMA_signal_3343), .B1_t (new_AGEMA_signal_3344), .B1_f (new_AGEMA_signal_3345), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3767), .Z1_t (new_AGEMA_signal_3768), .Z1_f (new_AGEMA_signal_3769) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3767), .B1_t (new_AGEMA_signal_3768), .B1_f (new_AGEMA_signal_3769), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4189), .Z1_t (new_AGEMA_signal_4190), .Z1_f (new_AGEMA_signal_4191) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4189), .A1_t (new_AGEMA_signal_4190), .A1_f (new_AGEMA_signal_4191), .B0_t (data_out_s0_t[50]), .B0_f (data_out_s0_f[50]), .B1_t (data_out_s1_t[50]), .B1_f (data_out_s1_f[50]), .Z0_t (data_out_s0_t[54]), .Z0_f (data_out_s0_f[54]), .Z1_t (data_out_s1_t[54]), .Z1_f (data_out_s1_f[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[51]), .A0_f (data_out_s0_f[51]), .A1_t (data_out_s1_t[51]), .A1_f (data_out_s1_f[51]), .B0_t (stateFF_inputPar[55]), .B0_f (new_AGEMA_signal_3346), .B1_t (new_AGEMA_signal_3347), .B1_f (new_AGEMA_signal_3348), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3770), .Z1_t (new_AGEMA_signal_3771), .Z1_f (new_AGEMA_signal_3772) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3770), .B1_t (new_AGEMA_signal_3771), .B1_f (new_AGEMA_signal_3772), .Z0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4192), .Z1_t (new_AGEMA_signal_4193), .Z1_f (new_AGEMA_signal_4194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4192), .A1_t (new_AGEMA_signal_4193), .A1_f (new_AGEMA_signal_4194), .B0_t (data_out_s0_t[51]), .B0_f (data_out_s0_f[51]), .B1_t (data_out_s1_t[51]), .B1_f (data_out_s1_f[51]), .Z0_t (data_out_s0_t[55]), .Z0_f (data_out_s0_f[55]), .Z1_t (data_out_s1_t[55]), .Z1_f (data_out_s1_f[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[52]), .A0_f (data_out_s0_f[52]), .A1_t (data_out_s1_t[52]), .A1_f (data_out_s1_f[52]), .B0_t (stateFF_inputPar[56]), .B0_f (new_AGEMA_signal_3349), .B1_t (new_AGEMA_signal_3350), .B1_f (new_AGEMA_signal_3351), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3773), .Z1_t (new_AGEMA_signal_3774), .Z1_f (new_AGEMA_signal_3775) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3773), .B1_t (new_AGEMA_signal_3774), .B1_f (new_AGEMA_signal_3775), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4195), .Z1_t (new_AGEMA_signal_4196), .Z1_f (new_AGEMA_signal_4197) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4195), .A1_t (new_AGEMA_signal_4196), .A1_f (new_AGEMA_signal_4197), .B0_t (data_out_s0_t[52]), .B0_f (data_out_s0_f[52]), .B1_t (data_out_s1_t[52]), .B1_f (data_out_s1_f[52]), .Z0_t (data_out_s0_t[56]), .Z0_f (data_out_s0_f[56]), .Z1_t (data_out_s1_t[56]), .Z1_f (data_out_s1_f[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[53]), .A0_f (data_out_s0_f[53]), .A1_t (data_out_s1_t[53]), .A1_f (data_out_s1_f[53]), .B0_t (stateFF_inputPar[57]), .B0_f (new_AGEMA_signal_3352), .B1_t (new_AGEMA_signal_3353), .B1_f (new_AGEMA_signal_3354), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3776), .Z1_t (new_AGEMA_signal_3777), .Z1_f (new_AGEMA_signal_3778) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3776), .B1_t (new_AGEMA_signal_3777), .B1_f (new_AGEMA_signal_3778), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4198), .Z1_t (new_AGEMA_signal_4199), .Z1_f (new_AGEMA_signal_4200) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4198), .A1_t (new_AGEMA_signal_4199), .A1_f (new_AGEMA_signal_4200), .B0_t (data_out_s0_t[53]), .B0_f (data_out_s0_f[53]), .B1_t (data_out_s1_t[53]), .B1_f (data_out_s1_f[53]), .Z0_t (data_out_s0_t[57]), .Z0_f (data_out_s0_f[57]), .Z1_t (data_out_s1_t[57]), .Z1_f (data_out_s1_f[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[54]), .A0_f (data_out_s0_f[54]), .A1_t (data_out_s1_t[54]), .A1_f (data_out_s1_f[54]), .B0_t (stateFF_inputPar[58]), .B0_f (new_AGEMA_signal_3355), .B1_t (new_AGEMA_signal_3356), .B1_f (new_AGEMA_signal_3357), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3779), .Z1_t (new_AGEMA_signal_3780), .Z1_f (new_AGEMA_signal_3781) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3779), .B1_t (new_AGEMA_signal_3780), .B1_f (new_AGEMA_signal_3781), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4201), .Z1_t (new_AGEMA_signal_4202), .Z1_f (new_AGEMA_signal_4203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4201), .A1_t (new_AGEMA_signal_4202), .A1_f (new_AGEMA_signal_4203), .B0_t (data_out_s0_t[54]), .B0_f (data_out_s0_f[54]), .B1_t (data_out_s1_t[54]), .B1_f (data_out_s1_f[54]), .Z0_t (data_out_s0_t[58]), .Z0_f (data_out_s0_f[58]), .Z1_t (data_out_s1_t[58]), .Z1_f (data_out_s1_f[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[55]), .A0_f (data_out_s0_f[55]), .A1_t (data_out_s1_t[55]), .A1_f (data_out_s1_f[55]), .B0_t (stateFF_inputPar[59]), .B0_f (new_AGEMA_signal_3358), .B1_t (new_AGEMA_signal_3359), .B1_f (new_AGEMA_signal_3360), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3782), .Z1_t (new_AGEMA_signal_3783), .Z1_f (new_AGEMA_signal_3784) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3782), .B1_t (new_AGEMA_signal_3783), .B1_f (new_AGEMA_signal_3784), .Z0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4204), .Z1_t (new_AGEMA_signal_4205), .Z1_f (new_AGEMA_signal_4206) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4204), .A1_t (new_AGEMA_signal_4205), .A1_f (new_AGEMA_signal_4206), .B0_t (data_out_s0_t[55]), .B0_f (data_out_s0_f[55]), .B1_t (data_out_s1_t[55]), .B1_f (data_out_s1_f[55]), .Z0_t (data_out_s0_t[59]), .Z0_f (data_out_s0_f[59]), .Z1_t (data_out_s1_t[59]), .Z1_f (data_out_s1_f[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[56]), .A0_f (data_out_s0_f[56]), .A1_t (data_out_s1_t[56]), .A1_f (data_out_s1_f[56]), .B0_t (stateFF_inputPar[60]), .B0_f (new_AGEMA_signal_3361), .B1_t (new_AGEMA_signal_3362), .B1_f (new_AGEMA_signal_3363), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3785), .Z1_t (new_AGEMA_signal_3786), .Z1_f (new_AGEMA_signal_3787) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3785), .B1_t (new_AGEMA_signal_3786), .B1_f (new_AGEMA_signal_3787), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4207), .Z1_t (new_AGEMA_signal_4208), .Z1_f (new_AGEMA_signal_4209) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4207), .A1_t (new_AGEMA_signal_4208), .A1_f (new_AGEMA_signal_4209), .B0_t (data_out_s0_t[56]), .B0_f (data_out_s0_f[56]), .B1_t (data_out_s1_t[56]), .B1_f (data_out_s1_f[56]), .Z0_t (data_out_s0_t[60]), .Z0_f (data_out_s0_f[60]), .Z1_t (data_out_s1_t[60]), .Z1_f (data_out_s1_f[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[57]), .A0_f (data_out_s0_f[57]), .A1_t (data_out_s1_t[57]), .A1_f (data_out_s1_f[57]), .B0_t (stateFF_inputPar[61]), .B0_f (new_AGEMA_signal_3364), .B1_t (new_AGEMA_signal_3365), .B1_f (new_AGEMA_signal_3366), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3788), .Z1_t (new_AGEMA_signal_3789), .Z1_f (new_AGEMA_signal_3790) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3788), .B1_t (new_AGEMA_signal_3789), .B1_f (new_AGEMA_signal_3790), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4210), .Z1_t (new_AGEMA_signal_4211), .Z1_f (new_AGEMA_signal_4212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4210), .A1_t (new_AGEMA_signal_4211), .A1_f (new_AGEMA_signal_4212), .B0_t (data_out_s0_t[57]), .B0_f (data_out_s0_f[57]), .B1_t (data_out_s1_t[57]), .B1_f (data_out_s1_f[57]), .Z0_t (data_out_s0_t[61]), .Z0_f (data_out_s0_f[61]), .Z1_t (data_out_s1_t[61]), .Z1_f (data_out_s1_f[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[58]), .A0_f (data_out_s0_f[58]), .A1_t (data_out_s1_t[58]), .A1_f (data_out_s1_f[58]), .B0_t (stateFF_inputPar[62]), .B0_f (new_AGEMA_signal_3367), .B1_t (new_AGEMA_signal_3368), .B1_f (new_AGEMA_signal_3369), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3791), .Z1_t (new_AGEMA_signal_3792), .Z1_f (new_AGEMA_signal_3793) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3791), .B1_t (new_AGEMA_signal_3792), .B1_f (new_AGEMA_signal_3793), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4213), .Z1_t (new_AGEMA_signal_4214), .Z1_f (new_AGEMA_signal_4215) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4213), .A1_t (new_AGEMA_signal_4214), .A1_f (new_AGEMA_signal_4215), .B0_t (data_out_s0_t[58]), .B0_f (data_out_s0_f[58]), .B1_t (data_out_s1_t[58]), .B1_f (data_out_s1_f[58]), .Z0_t (data_out_s0_t[62]), .Z0_f (data_out_s0_f[62]), .Z1_t (data_out_s1_t[62]), .Z1_f (data_out_s1_f[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[59]), .A0_f (data_out_s0_f[59]), .A1_t (data_out_s1_t[59]), .A1_f (data_out_s1_f[59]), .B0_t (stateFF_inputPar[63]), .B0_f (new_AGEMA_signal_3370), .B1_t (new_AGEMA_signal_3371), .B1_f (new_AGEMA_signal_3372), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3794), .Z1_t (new_AGEMA_signal_3795), .Z1_f (new_AGEMA_signal_3796) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3794), .B1_t (new_AGEMA_signal_3795), .B1_f (new_AGEMA_signal_3796), .Z0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4216), .Z1_t (new_AGEMA_signal_4217), .Z1_f (new_AGEMA_signal_4218) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4216), .A1_t (new_AGEMA_signal_4217), .A1_f (new_AGEMA_signal_4218), .B0_t (data_out_s0_t[59]), .B0_f (data_out_s0_f[59]), .B1_t (data_out_s1_t[59]), .B1_f (data_out_s1_f[59]), .Z0_t (data_out_s0_t[63]), .Z0_f (data_out_s0_f[63]), .Z1_t (data_out_s1_t[63]), .Z1_f (data_out_s1_f[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_XOR1_U1 ( .A0_t (data_out_s0_t[0]), .A0_f (data_out_s0_f[0]), .A1_t (data_out_s1_t[0]), .A1_f (data_out_s1_f[0]), .B0_t (data_in_s0_t[0]), .B0_f (data_in_s0_f[0]), .B1_t (data_in_s1_t[0]), .B1_f (data_in_s1_f[0]), .Z0_t (stateFF_MUX_inputPar_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_1496), .Z1_t (new_AGEMA_signal_1497), .Z1_f (new_AGEMA_signal_1498) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_1496), .B1_t (new_AGEMA_signal_1497), .B1_f (new_AGEMA_signal_1498), .Z0_t (stateFF_MUX_inputPar_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_2721), .Z1_t (new_AGEMA_signal_2722), .Z1_f (new_AGEMA_signal_2723) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_0_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_2721), .A1_t (new_AGEMA_signal_2722), .A1_f (new_AGEMA_signal_2723), .B0_t (data_out_s0_t[0]), .B0_f (data_out_s0_f[0]), .B1_t (data_out_s1_t[0]), .B1_f (data_out_s1_f[0]), .Z0_t (stateFF_inputPar[0]), .Z0_f (new_AGEMA_signal_3181), .Z1_t (new_AGEMA_signal_3182), .Z1_f (new_AGEMA_signal_3183) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_XOR1_U1 ( .A0_t (data_out_s0_t[4]), .A0_f (data_out_s0_f[4]), .A1_t (data_out_s1_t[4]), .A1_f (data_out_s1_f[4]), .B0_t (data_in_s0_t[1]), .B0_f (data_in_s0_f[1]), .B1_t (data_in_s1_t[1]), .B1_f (data_in_s1_f[1]), .Z0_t (stateFF_MUX_inputPar_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_1505), .Z1_t (new_AGEMA_signal_1506), .Z1_f (new_AGEMA_signal_1507) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_1505), .B1_t (new_AGEMA_signal_1506), .B1_f (new_AGEMA_signal_1507), .Z0_t (stateFF_MUX_inputPar_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_2724), .Z1_t (new_AGEMA_signal_2725), .Z1_f (new_AGEMA_signal_2726) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_1_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_2724), .A1_t (new_AGEMA_signal_2725), .A1_f (new_AGEMA_signal_2726), .B0_t (data_out_s0_t[4]), .B0_f (data_out_s0_f[4]), .B1_t (data_out_s1_t[4]), .B1_f (data_out_s1_f[4]), .Z0_t (stateFF_inputPar[1]), .Z0_f (new_AGEMA_signal_3184), .Z1_t (new_AGEMA_signal_3185), .Z1_f (new_AGEMA_signal_3186) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_XOR1_U1 ( .A0_t (data_out_s0_t[8]), .A0_f (data_out_s0_f[8]), .A1_t (data_out_s1_t[8]), .A1_f (data_out_s1_f[8]), .B0_t (data_in_s0_t[2]), .B0_f (data_in_s0_f[2]), .B1_t (data_in_s1_t[2]), .B1_f (data_in_s1_f[2]), .Z0_t (stateFF_MUX_inputPar_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_1514), .Z1_t (new_AGEMA_signal_1515), .Z1_f (new_AGEMA_signal_1516) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_1514), .B1_t (new_AGEMA_signal_1515), .B1_f (new_AGEMA_signal_1516), .Z0_t (stateFF_MUX_inputPar_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_2727), .Z1_t (new_AGEMA_signal_2728), .Z1_f (new_AGEMA_signal_2729) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_2_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_2727), .A1_t (new_AGEMA_signal_2728), .A1_f (new_AGEMA_signal_2729), .B0_t (data_out_s0_t[8]), .B0_f (data_out_s0_f[8]), .B1_t (data_out_s1_t[8]), .B1_f (data_out_s1_f[8]), .Z0_t (stateFF_inputPar[2]), .Z0_f (new_AGEMA_signal_3187), .Z1_t (new_AGEMA_signal_3188), .Z1_f (new_AGEMA_signal_3189) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_XOR1_U1 ( .A0_t (data_out_s0_t[12]), .A0_f (data_out_s0_f[12]), .A1_t (data_out_s1_t[12]), .A1_f (data_out_s1_f[12]), .B0_t (data_in_s0_t[3]), .B0_f (data_in_s0_f[3]), .B1_t (data_in_s1_t[3]), .B1_f (data_in_s1_f[3]), .Z0_t (stateFF_MUX_inputPar_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_1523), .Z1_t (new_AGEMA_signal_1524), .Z1_f (new_AGEMA_signal_1525) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_1523), .B1_t (new_AGEMA_signal_1524), .B1_f (new_AGEMA_signal_1525), .Z0_t (stateFF_MUX_inputPar_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_2730), .Z1_t (new_AGEMA_signal_2731), .Z1_f (new_AGEMA_signal_2732) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_3_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_2730), .A1_t (new_AGEMA_signal_2731), .A1_f (new_AGEMA_signal_2732), .B0_t (data_out_s0_t[12]), .B0_f (data_out_s0_f[12]), .B1_t (data_out_s1_t[12]), .B1_f (data_out_s1_f[12]), .Z0_t (stateFF_inputPar[3]), .Z0_f (new_AGEMA_signal_3190), .Z1_t (new_AGEMA_signal_3191), .Z1_f (new_AGEMA_signal_3192) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_XOR1_U1 ( .A0_t (data_out_s0_t[16]), .A0_f (data_out_s0_f[16]), .A1_t (data_out_s1_t[16]), .A1_f (data_out_s1_f[16]), .B0_t (data_in_s0_t[4]), .B0_f (data_in_s0_f[4]), .B1_t (data_in_s1_t[4]), .B1_f (data_in_s1_f[4]), .Z0_t (stateFF_MUX_inputPar_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_1532), .Z1_t (new_AGEMA_signal_1533), .Z1_f (new_AGEMA_signal_1534) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_1532), .B1_t (new_AGEMA_signal_1533), .B1_f (new_AGEMA_signal_1534), .Z0_t (stateFF_MUX_inputPar_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_2733), .Z1_t (new_AGEMA_signal_2734), .Z1_f (new_AGEMA_signal_2735) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_4_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_2733), .A1_t (new_AGEMA_signal_2734), .A1_f (new_AGEMA_signal_2735), .B0_t (data_out_s0_t[16]), .B0_f (data_out_s0_f[16]), .B1_t (data_out_s1_t[16]), .B1_f (data_out_s1_f[16]), .Z0_t (stateFF_inputPar[4]), .Z0_f (new_AGEMA_signal_3193), .Z1_t (new_AGEMA_signal_3194), .Z1_f (new_AGEMA_signal_3195) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_XOR1_U1 ( .A0_t (data_out_s0_t[20]), .A0_f (data_out_s0_f[20]), .A1_t (data_out_s1_t[20]), .A1_f (data_out_s1_f[20]), .B0_t (data_in_s0_t[5]), .B0_f (data_in_s0_f[5]), .B1_t (data_in_s1_t[5]), .B1_f (data_in_s1_f[5]), .Z0_t (stateFF_MUX_inputPar_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_1541), .Z1_t (new_AGEMA_signal_1542), .Z1_f (new_AGEMA_signal_1543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_1541), .B1_t (new_AGEMA_signal_1542), .B1_f (new_AGEMA_signal_1543), .Z0_t (stateFF_MUX_inputPar_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_2736), .Z1_t (new_AGEMA_signal_2737), .Z1_f (new_AGEMA_signal_2738) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_5_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_2736), .A1_t (new_AGEMA_signal_2737), .A1_f (new_AGEMA_signal_2738), .B0_t (data_out_s0_t[20]), .B0_f (data_out_s0_f[20]), .B1_t (data_out_s1_t[20]), .B1_f (data_out_s1_f[20]), .Z0_t (stateFF_inputPar[5]), .Z0_f (new_AGEMA_signal_3196), .Z1_t (new_AGEMA_signal_3197), .Z1_f (new_AGEMA_signal_3198) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_XOR1_U1 ( .A0_t (data_out_s0_t[24]), .A0_f (data_out_s0_f[24]), .A1_t (data_out_s1_t[24]), .A1_f (data_out_s1_f[24]), .B0_t (data_in_s0_t[6]), .B0_f (data_in_s0_f[6]), .B1_t (data_in_s1_t[6]), .B1_f (data_in_s1_f[6]), .Z0_t (stateFF_MUX_inputPar_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_1550), .Z1_t (new_AGEMA_signal_1551), .Z1_f (new_AGEMA_signal_1552) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_1550), .B1_t (new_AGEMA_signal_1551), .B1_f (new_AGEMA_signal_1552), .Z0_t (stateFF_MUX_inputPar_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_2739), .Z1_t (new_AGEMA_signal_2740), .Z1_f (new_AGEMA_signal_2741) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_6_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_2739), .A1_t (new_AGEMA_signal_2740), .A1_f (new_AGEMA_signal_2741), .B0_t (data_out_s0_t[24]), .B0_f (data_out_s0_f[24]), .B1_t (data_out_s1_t[24]), .B1_f (data_out_s1_f[24]), .Z0_t (stateFF_inputPar[6]), .Z0_f (new_AGEMA_signal_3199), .Z1_t (new_AGEMA_signal_3200), .Z1_f (new_AGEMA_signal_3201) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_XOR1_U1 ( .A0_t (data_out_s0_t[28]), .A0_f (data_out_s0_f[28]), .A1_t (data_out_s1_t[28]), .A1_f (data_out_s1_f[28]), .B0_t (data_in_s0_t[7]), .B0_f (data_in_s0_f[7]), .B1_t (data_in_s1_t[7]), .B1_f (data_in_s1_f[7]), .Z0_t (stateFF_MUX_inputPar_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_1559), .Z1_t (new_AGEMA_signal_1560), .Z1_f (new_AGEMA_signal_1561) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_1559), .B1_t (new_AGEMA_signal_1560), .B1_f (new_AGEMA_signal_1561), .Z0_t (stateFF_MUX_inputPar_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_2742), .Z1_t (new_AGEMA_signal_2743), .Z1_f (new_AGEMA_signal_2744) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_7_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_2742), .A1_t (new_AGEMA_signal_2743), .A1_f (new_AGEMA_signal_2744), .B0_t (data_out_s0_t[28]), .B0_f (data_out_s0_f[28]), .B1_t (data_out_s1_t[28]), .B1_f (data_out_s1_f[28]), .Z0_t (stateFF_inputPar[7]), .Z0_f (new_AGEMA_signal_3202), .Z1_t (new_AGEMA_signal_3203), .Z1_f (new_AGEMA_signal_3204) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_XOR1_U1 ( .A0_t (data_out_s0_t[32]), .A0_f (data_out_s0_f[32]), .A1_t (data_out_s1_t[32]), .A1_f (data_out_s1_f[32]), .B0_t (data_in_s0_t[8]), .B0_f (data_in_s0_f[8]), .B1_t (data_in_s1_t[8]), .B1_f (data_in_s1_f[8]), .Z0_t (stateFF_MUX_inputPar_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_1568), .Z1_t (new_AGEMA_signal_1569), .Z1_f (new_AGEMA_signal_1570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_1568), .B1_t (new_AGEMA_signal_1569), .B1_f (new_AGEMA_signal_1570), .Z0_t (stateFF_MUX_inputPar_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_2745), .Z1_t (new_AGEMA_signal_2746), .Z1_f (new_AGEMA_signal_2747) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_8_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_2745), .A1_t (new_AGEMA_signal_2746), .A1_f (new_AGEMA_signal_2747), .B0_t (data_out_s0_t[32]), .B0_f (data_out_s0_f[32]), .B1_t (data_out_s1_t[32]), .B1_f (data_out_s1_f[32]), .Z0_t (stateFF_inputPar[8]), .Z0_f (new_AGEMA_signal_3205), .Z1_t (new_AGEMA_signal_3206), .Z1_f (new_AGEMA_signal_3207) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_XOR1_U1 ( .A0_t (data_out_s0_t[36]), .A0_f (data_out_s0_f[36]), .A1_t (data_out_s1_t[36]), .A1_f (data_out_s1_f[36]), .B0_t (data_in_s0_t[9]), .B0_f (data_in_s0_f[9]), .B1_t (data_in_s1_t[9]), .B1_f (data_in_s1_f[9]), .Z0_t (stateFF_MUX_inputPar_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_1577), .Z1_t (new_AGEMA_signal_1578), .Z1_f (new_AGEMA_signal_1579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_1577), .B1_t (new_AGEMA_signal_1578), .B1_f (new_AGEMA_signal_1579), .Z0_t (stateFF_MUX_inputPar_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_2748), .Z1_t (new_AGEMA_signal_2749), .Z1_f (new_AGEMA_signal_2750) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_9_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_2748), .A1_t (new_AGEMA_signal_2749), .A1_f (new_AGEMA_signal_2750), .B0_t (data_out_s0_t[36]), .B0_f (data_out_s0_f[36]), .B1_t (data_out_s1_t[36]), .B1_f (data_out_s1_f[36]), .Z0_t (stateFF_inputPar[9]), .Z0_f (new_AGEMA_signal_3208), .Z1_t (new_AGEMA_signal_3209), .Z1_f (new_AGEMA_signal_3210) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_XOR1_U1 ( .A0_t (data_out_s0_t[40]), .A0_f (data_out_s0_f[40]), .A1_t (data_out_s1_t[40]), .A1_f (data_out_s1_f[40]), .B0_t (data_in_s0_t[10]), .B0_f (data_in_s0_f[10]), .B1_t (data_in_s1_t[10]), .B1_f (data_in_s1_f[10]), .Z0_t (stateFF_MUX_inputPar_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_1586), .Z1_t (new_AGEMA_signal_1587), .Z1_f (new_AGEMA_signal_1588) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_1586), .B1_t (new_AGEMA_signal_1587), .B1_f (new_AGEMA_signal_1588), .Z0_t (stateFF_MUX_inputPar_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_2751), .Z1_t (new_AGEMA_signal_2752), .Z1_f (new_AGEMA_signal_2753) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_10_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_2751), .A1_t (new_AGEMA_signal_2752), .A1_f (new_AGEMA_signal_2753), .B0_t (data_out_s0_t[40]), .B0_f (data_out_s0_f[40]), .B1_t (data_out_s1_t[40]), .B1_f (data_out_s1_f[40]), .Z0_t (stateFF_inputPar[10]), .Z0_f (new_AGEMA_signal_3211), .Z1_t (new_AGEMA_signal_3212), .Z1_f (new_AGEMA_signal_3213) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_XOR1_U1 ( .A0_t (data_out_s0_t[44]), .A0_f (data_out_s0_f[44]), .A1_t (data_out_s1_t[44]), .A1_f (data_out_s1_f[44]), .B0_t (data_in_s0_t[11]), .B0_f (data_in_s0_f[11]), .B1_t (data_in_s1_t[11]), .B1_f (data_in_s1_f[11]), .Z0_t (stateFF_MUX_inputPar_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_1595), .Z1_t (new_AGEMA_signal_1596), .Z1_f (new_AGEMA_signal_1597) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_1595), .B1_t (new_AGEMA_signal_1596), .B1_f (new_AGEMA_signal_1597), .Z0_t (stateFF_MUX_inputPar_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_2754), .Z1_t (new_AGEMA_signal_2755), .Z1_f (new_AGEMA_signal_2756) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_11_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_2754), .A1_t (new_AGEMA_signal_2755), .A1_f (new_AGEMA_signal_2756), .B0_t (data_out_s0_t[44]), .B0_f (data_out_s0_f[44]), .B1_t (data_out_s1_t[44]), .B1_f (data_out_s1_f[44]), .Z0_t (stateFF_inputPar[11]), .Z0_f (new_AGEMA_signal_3214), .Z1_t (new_AGEMA_signal_3215), .Z1_f (new_AGEMA_signal_3216) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_XOR1_U1 ( .A0_t (data_out_s0_t[48]), .A0_f (data_out_s0_f[48]), .A1_t (data_out_s1_t[48]), .A1_f (data_out_s1_f[48]), .B0_t (data_in_s0_t[12]), .B0_f (data_in_s0_f[12]), .B1_t (data_in_s1_t[12]), .B1_f (data_in_s1_f[12]), .Z0_t (stateFF_MUX_inputPar_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_1604), .Z1_t (new_AGEMA_signal_1605), .Z1_f (new_AGEMA_signal_1606) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_1604), .B1_t (new_AGEMA_signal_1605), .B1_f (new_AGEMA_signal_1606), .Z0_t (stateFF_MUX_inputPar_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_2757), .Z1_t (new_AGEMA_signal_2758), .Z1_f (new_AGEMA_signal_2759) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_12_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_2757), .A1_t (new_AGEMA_signal_2758), .A1_f (new_AGEMA_signal_2759), .B0_t (data_out_s0_t[48]), .B0_f (data_out_s0_f[48]), .B1_t (data_out_s1_t[48]), .B1_f (data_out_s1_f[48]), .Z0_t (stateFF_inputPar[12]), .Z0_f (new_AGEMA_signal_3217), .Z1_t (new_AGEMA_signal_3218), .Z1_f (new_AGEMA_signal_3219) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_XOR1_U1 ( .A0_t (data_out_s0_t[52]), .A0_f (data_out_s0_f[52]), .A1_t (data_out_s1_t[52]), .A1_f (data_out_s1_f[52]), .B0_t (data_in_s0_t[13]), .B0_f (data_in_s0_f[13]), .B1_t (data_in_s1_t[13]), .B1_f (data_in_s1_f[13]), .Z0_t (stateFF_MUX_inputPar_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_1613), .Z1_t (new_AGEMA_signal_1614), .Z1_f (new_AGEMA_signal_1615) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_1613), .B1_t (new_AGEMA_signal_1614), .B1_f (new_AGEMA_signal_1615), .Z0_t (stateFF_MUX_inputPar_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_2760), .Z1_t (new_AGEMA_signal_2761), .Z1_f (new_AGEMA_signal_2762) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_13_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_2760), .A1_t (new_AGEMA_signal_2761), .A1_f (new_AGEMA_signal_2762), .B0_t (data_out_s0_t[52]), .B0_f (data_out_s0_f[52]), .B1_t (data_out_s1_t[52]), .B1_f (data_out_s1_f[52]), .Z0_t (stateFF_inputPar[13]), .Z0_f (new_AGEMA_signal_3220), .Z1_t (new_AGEMA_signal_3221), .Z1_f (new_AGEMA_signal_3222) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_XOR1_U1 ( .A0_t (data_out_s0_t[56]), .A0_f (data_out_s0_f[56]), .A1_t (data_out_s1_t[56]), .A1_f (data_out_s1_f[56]), .B0_t (data_in_s0_t[14]), .B0_f (data_in_s0_f[14]), .B1_t (data_in_s1_t[14]), .B1_f (data_in_s1_f[14]), .Z0_t (stateFF_MUX_inputPar_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_1622), .Z1_t (new_AGEMA_signal_1623), .Z1_f (new_AGEMA_signal_1624) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_1622), .B1_t (new_AGEMA_signal_1623), .B1_f (new_AGEMA_signal_1624), .Z0_t (stateFF_MUX_inputPar_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_2763), .Z1_t (new_AGEMA_signal_2764), .Z1_f (new_AGEMA_signal_2765) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_14_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_2763), .A1_t (new_AGEMA_signal_2764), .A1_f (new_AGEMA_signal_2765), .B0_t (data_out_s0_t[56]), .B0_f (data_out_s0_f[56]), .B1_t (data_out_s1_t[56]), .B1_f (data_out_s1_f[56]), .Z0_t (stateFF_inputPar[14]), .Z0_f (new_AGEMA_signal_3223), .Z1_t (new_AGEMA_signal_3224), .Z1_f (new_AGEMA_signal_3225) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_XOR1_U1 ( .A0_t (data_out_s0_t[60]), .A0_f (data_out_s0_f[60]), .A1_t (data_out_s1_t[60]), .A1_f (data_out_s1_f[60]), .B0_t (data_in_s0_t[15]), .B0_f (data_in_s0_f[15]), .B1_t (data_in_s1_t[15]), .B1_f (data_in_s1_f[15]), .Z0_t (stateFF_MUX_inputPar_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_1628), .Z1_t (new_AGEMA_signal_1629), .Z1_f (new_AGEMA_signal_1630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_1628), .B1_t (new_AGEMA_signal_1629), .B1_f (new_AGEMA_signal_1630), .Z0_t (stateFF_MUX_inputPar_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_2766), .Z1_t (new_AGEMA_signal_2767), .Z1_f (new_AGEMA_signal_2768) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_15_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_2766), .A1_t (new_AGEMA_signal_2767), .A1_f (new_AGEMA_signal_2768), .B0_t (data_out_s0_t[60]), .B0_f (data_out_s0_f[60]), .B1_t (data_out_s1_t[60]), .B1_f (data_out_s1_f[60]), .Z0_t (stateFF_inputPar[15]), .Z0_f (new_AGEMA_signal_3226), .Z1_t (new_AGEMA_signal_3227), .Z1_f (new_AGEMA_signal_3228) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_XOR1_U1 ( .A0_t (data_out_s0_t[1]), .A0_f (data_out_s0_f[1]), .A1_t (data_out_s1_t[1]), .A1_f (data_out_s1_f[1]), .B0_t (data_in_s0_t[16]), .B0_f (data_in_s0_f[16]), .B1_t (data_in_s1_t[16]), .B1_f (data_in_s1_f[16]), .Z0_t (stateFF_MUX_inputPar_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_1637), .Z1_t (new_AGEMA_signal_1638), .Z1_f (new_AGEMA_signal_1639) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_1637), .B1_t (new_AGEMA_signal_1638), .B1_f (new_AGEMA_signal_1639), .Z0_t (stateFF_MUX_inputPar_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_2769), .Z1_t (new_AGEMA_signal_2770), .Z1_f (new_AGEMA_signal_2771) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_16_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_2769), .A1_t (new_AGEMA_signal_2770), .A1_f (new_AGEMA_signal_2771), .B0_t (data_out_s0_t[1]), .B0_f (data_out_s0_f[1]), .B1_t (data_out_s1_t[1]), .B1_f (data_out_s1_f[1]), .Z0_t (stateFF_inputPar[16]), .Z0_f (new_AGEMA_signal_3229), .Z1_t (new_AGEMA_signal_3230), .Z1_f (new_AGEMA_signal_3231) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_XOR1_U1 ( .A0_t (data_out_s0_t[5]), .A0_f (data_out_s0_f[5]), .A1_t (data_out_s1_t[5]), .A1_f (data_out_s1_f[5]), .B0_t (data_in_s0_t[17]), .B0_f (data_in_s0_f[17]), .B1_t (data_in_s1_t[17]), .B1_f (data_in_s1_f[17]), .Z0_t (stateFF_MUX_inputPar_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_1646), .Z1_t (new_AGEMA_signal_1647), .Z1_f (new_AGEMA_signal_1648) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_1646), .B1_t (new_AGEMA_signal_1647), .B1_f (new_AGEMA_signal_1648), .Z0_t (stateFF_MUX_inputPar_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_2772), .Z1_t (new_AGEMA_signal_2773), .Z1_f (new_AGEMA_signal_2774) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_17_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_2772), .A1_t (new_AGEMA_signal_2773), .A1_f (new_AGEMA_signal_2774), .B0_t (data_out_s0_t[5]), .B0_f (data_out_s0_f[5]), .B1_t (data_out_s1_t[5]), .B1_f (data_out_s1_f[5]), .Z0_t (stateFF_inputPar[17]), .Z0_f (new_AGEMA_signal_3232), .Z1_t (new_AGEMA_signal_3233), .Z1_f (new_AGEMA_signal_3234) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_XOR1_U1 ( .A0_t (data_out_s0_t[9]), .A0_f (data_out_s0_f[9]), .A1_t (data_out_s1_t[9]), .A1_f (data_out_s1_f[9]), .B0_t (data_in_s0_t[18]), .B0_f (data_in_s0_f[18]), .B1_t (data_in_s1_t[18]), .B1_f (data_in_s1_f[18]), .Z0_t (stateFF_MUX_inputPar_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_1655), .Z1_t (new_AGEMA_signal_1656), .Z1_f (new_AGEMA_signal_1657) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_1655), .B1_t (new_AGEMA_signal_1656), .B1_f (new_AGEMA_signal_1657), .Z0_t (stateFF_MUX_inputPar_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_2775), .Z1_t (new_AGEMA_signal_2776), .Z1_f (new_AGEMA_signal_2777) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_18_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_2775), .A1_t (new_AGEMA_signal_2776), .A1_f (new_AGEMA_signal_2777), .B0_t (data_out_s0_t[9]), .B0_f (data_out_s0_f[9]), .B1_t (data_out_s1_t[9]), .B1_f (data_out_s1_f[9]), .Z0_t (stateFF_inputPar[18]), .Z0_f (new_AGEMA_signal_3235), .Z1_t (new_AGEMA_signal_3236), .Z1_f (new_AGEMA_signal_3237) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_XOR1_U1 ( .A0_t (data_out_s0_t[13]), .A0_f (data_out_s0_f[13]), .A1_t (data_out_s1_t[13]), .A1_f (data_out_s1_f[13]), .B0_t (data_in_s0_t[19]), .B0_f (data_in_s0_f[19]), .B1_t (data_in_s1_t[19]), .B1_f (data_in_s1_f[19]), .Z0_t (stateFF_MUX_inputPar_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_1664), .Z1_t (new_AGEMA_signal_1665), .Z1_f (new_AGEMA_signal_1666) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_1664), .B1_t (new_AGEMA_signal_1665), .B1_f (new_AGEMA_signal_1666), .Z0_t (stateFF_MUX_inputPar_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_2778), .Z1_t (new_AGEMA_signal_2779), .Z1_f (new_AGEMA_signal_2780) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_19_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_2778), .A1_t (new_AGEMA_signal_2779), .A1_f (new_AGEMA_signal_2780), .B0_t (data_out_s0_t[13]), .B0_f (data_out_s0_f[13]), .B1_t (data_out_s1_t[13]), .B1_f (data_out_s1_f[13]), .Z0_t (stateFF_inputPar[19]), .Z0_f (new_AGEMA_signal_3238), .Z1_t (new_AGEMA_signal_3239), .Z1_f (new_AGEMA_signal_3240) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_XOR1_U1 ( .A0_t (data_out_s0_t[17]), .A0_f (data_out_s0_f[17]), .A1_t (data_out_s1_t[17]), .A1_f (data_out_s1_f[17]), .B0_t (data_in_s0_t[20]), .B0_f (data_in_s0_f[20]), .B1_t (data_in_s1_t[20]), .B1_f (data_in_s1_f[20]), .Z0_t (stateFF_MUX_inputPar_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_1673), .Z1_t (new_AGEMA_signal_1674), .Z1_f (new_AGEMA_signal_1675) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_1673), .B1_t (new_AGEMA_signal_1674), .B1_f (new_AGEMA_signal_1675), .Z0_t (stateFF_MUX_inputPar_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_2781), .Z1_t (new_AGEMA_signal_2782), .Z1_f (new_AGEMA_signal_2783) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_20_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_2781), .A1_t (new_AGEMA_signal_2782), .A1_f (new_AGEMA_signal_2783), .B0_t (data_out_s0_t[17]), .B0_f (data_out_s0_f[17]), .B1_t (data_out_s1_t[17]), .B1_f (data_out_s1_f[17]), .Z0_t (stateFF_inputPar[20]), .Z0_f (new_AGEMA_signal_3241), .Z1_t (new_AGEMA_signal_3242), .Z1_f (new_AGEMA_signal_3243) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_XOR1_U1 ( .A0_t (data_out_s0_t[21]), .A0_f (data_out_s0_f[21]), .A1_t (data_out_s1_t[21]), .A1_f (data_out_s1_f[21]), .B0_t (data_in_s0_t[21]), .B0_f (data_in_s0_f[21]), .B1_t (data_in_s1_t[21]), .B1_f (data_in_s1_f[21]), .Z0_t (stateFF_MUX_inputPar_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_1682), .Z1_t (new_AGEMA_signal_1683), .Z1_f (new_AGEMA_signal_1684) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_1682), .B1_t (new_AGEMA_signal_1683), .B1_f (new_AGEMA_signal_1684), .Z0_t (stateFF_MUX_inputPar_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_2784), .Z1_t (new_AGEMA_signal_2785), .Z1_f (new_AGEMA_signal_2786) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_21_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_2784), .A1_t (new_AGEMA_signal_2785), .A1_f (new_AGEMA_signal_2786), .B0_t (data_out_s0_t[21]), .B0_f (data_out_s0_f[21]), .B1_t (data_out_s1_t[21]), .B1_f (data_out_s1_f[21]), .Z0_t (stateFF_inputPar[21]), .Z0_f (new_AGEMA_signal_3244), .Z1_t (new_AGEMA_signal_3245), .Z1_f (new_AGEMA_signal_3246) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_XOR1_U1 ( .A0_t (data_out_s0_t[25]), .A0_f (data_out_s0_f[25]), .A1_t (data_out_s1_t[25]), .A1_f (data_out_s1_f[25]), .B0_t (data_in_s0_t[22]), .B0_f (data_in_s0_f[22]), .B1_t (data_in_s1_t[22]), .B1_f (data_in_s1_f[22]), .Z0_t (stateFF_MUX_inputPar_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_1691), .Z1_t (new_AGEMA_signal_1692), .Z1_f (new_AGEMA_signal_1693) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_1691), .B1_t (new_AGEMA_signal_1692), .B1_f (new_AGEMA_signal_1693), .Z0_t (stateFF_MUX_inputPar_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_2787), .Z1_t (new_AGEMA_signal_2788), .Z1_f (new_AGEMA_signal_2789) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_22_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_2787), .A1_t (new_AGEMA_signal_2788), .A1_f (new_AGEMA_signal_2789), .B0_t (data_out_s0_t[25]), .B0_f (data_out_s0_f[25]), .B1_t (data_out_s1_t[25]), .B1_f (data_out_s1_f[25]), .Z0_t (stateFF_inputPar[22]), .Z0_f (new_AGEMA_signal_3247), .Z1_t (new_AGEMA_signal_3248), .Z1_f (new_AGEMA_signal_3249) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_XOR1_U1 ( .A0_t (data_out_s0_t[29]), .A0_f (data_out_s0_f[29]), .A1_t (data_out_s1_t[29]), .A1_f (data_out_s1_f[29]), .B0_t (data_in_s0_t[23]), .B0_f (data_in_s0_f[23]), .B1_t (data_in_s1_t[23]), .B1_f (data_in_s1_f[23]), .Z0_t (stateFF_MUX_inputPar_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_1700), .Z1_t (new_AGEMA_signal_1701), .Z1_f (new_AGEMA_signal_1702) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_1700), .B1_t (new_AGEMA_signal_1701), .B1_f (new_AGEMA_signal_1702), .Z0_t (stateFF_MUX_inputPar_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_2790), .Z1_t (new_AGEMA_signal_2791), .Z1_f (new_AGEMA_signal_2792) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_23_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_2790), .A1_t (new_AGEMA_signal_2791), .A1_f (new_AGEMA_signal_2792), .B0_t (data_out_s0_t[29]), .B0_f (data_out_s0_f[29]), .B1_t (data_out_s1_t[29]), .B1_f (data_out_s1_f[29]), .Z0_t (stateFF_inputPar[23]), .Z0_f (new_AGEMA_signal_3250), .Z1_t (new_AGEMA_signal_3251), .Z1_f (new_AGEMA_signal_3252) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_XOR1_U1 ( .A0_t (data_out_s0_t[33]), .A0_f (data_out_s0_f[33]), .A1_t (data_out_s1_t[33]), .A1_f (data_out_s1_f[33]), .B0_t (data_in_s0_t[24]), .B0_f (data_in_s0_f[24]), .B1_t (data_in_s1_t[24]), .B1_f (data_in_s1_f[24]), .Z0_t (stateFF_MUX_inputPar_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_1709), .Z1_t (new_AGEMA_signal_1710), .Z1_f (new_AGEMA_signal_1711) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_1709), .B1_t (new_AGEMA_signal_1710), .B1_f (new_AGEMA_signal_1711), .Z0_t (stateFF_MUX_inputPar_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_2793), .Z1_t (new_AGEMA_signal_2794), .Z1_f (new_AGEMA_signal_2795) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_24_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_2793), .A1_t (new_AGEMA_signal_2794), .A1_f (new_AGEMA_signal_2795), .B0_t (data_out_s0_t[33]), .B0_f (data_out_s0_f[33]), .B1_t (data_out_s1_t[33]), .B1_f (data_out_s1_f[33]), .Z0_t (stateFF_inputPar[24]), .Z0_f (new_AGEMA_signal_3253), .Z1_t (new_AGEMA_signal_3254), .Z1_f (new_AGEMA_signal_3255) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_XOR1_U1 ( .A0_t (data_out_s0_t[37]), .A0_f (data_out_s0_f[37]), .A1_t (data_out_s1_t[37]), .A1_f (data_out_s1_f[37]), .B0_t (data_in_s0_t[25]), .B0_f (data_in_s0_f[25]), .B1_t (data_in_s1_t[25]), .B1_f (data_in_s1_f[25]), .Z0_t (stateFF_MUX_inputPar_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_1718), .Z1_t (new_AGEMA_signal_1719), .Z1_f (new_AGEMA_signal_1720) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_1718), .B1_t (new_AGEMA_signal_1719), .B1_f (new_AGEMA_signal_1720), .Z0_t (stateFF_MUX_inputPar_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_2796), .Z1_t (new_AGEMA_signal_2797), .Z1_f (new_AGEMA_signal_2798) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_25_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_2796), .A1_t (new_AGEMA_signal_2797), .A1_f (new_AGEMA_signal_2798), .B0_t (data_out_s0_t[37]), .B0_f (data_out_s0_f[37]), .B1_t (data_out_s1_t[37]), .B1_f (data_out_s1_f[37]), .Z0_t (stateFF_inputPar[25]), .Z0_f (new_AGEMA_signal_3256), .Z1_t (new_AGEMA_signal_3257), .Z1_f (new_AGEMA_signal_3258) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_XOR1_U1 ( .A0_t (data_out_s0_t[41]), .A0_f (data_out_s0_f[41]), .A1_t (data_out_s1_t[41]), .A1_f (data_out_s1_f[41]), .B0_t (data_in_s0_t[26]), .B0_f (data_in_s0_f[26]), .B1_t (data_in_s1_t[26]), .B1_f (data_in_s1_f[26]), .Z0_t (stateFF_MUX_inputPar_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_1727), .Z1_t (new_AGEMA_signal_1728), .Z1_f (new_AGEMA_signal_1729) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_1727), .B1_t (new_AGEMA_signal_1728), .B1_f (new_AGEMA_signal_1729), .Z0_t (stateFF_MUX_inputPar_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_2799), .Z1_t (new_AGEMA_signal_2800), .Z1_f (new_AGEMA_signal_2801) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_26_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_2799), .A1_t (new_AGEMA_signal_2800), .A1_f (new_AGEMA_signal_2801), .B0_t (data_out_s0_t[41]), .B0_f (data_out_s0_f[41]), .B1_t (data_out_s1_t[41]), .B1_f (data_out_s1_f[41]), .Z0_t (stateFF_inputPar[26]), .Z0_f (new_AGEMA_signal_3259), .Z1_t (new_AGEMA_signal_3260), .Z1_f (new_AGEMA_signal_3261) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_XOR1_U1 ( .A0_t (data_out_s0_t[45]), .A0_f (data_out_s0_f[45]), .A1_t (data_out_s1_t[45]), .A1_f (data_out_s1_f[45]), .B0_t (data_in_s0_t[27]), .B0_f (data_in_s0_f[27]), .B1_t (data_in_s1_t[27]), .B1_f (data_in_s1_f[27]), .Z0_t (stateFF_MUX_inputPar_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_1736), .Z1_t (new_AGEMA_signal_1737), .Z1_f (new_AGEMA_signal_1738) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_1736), .B1_t (new_AGEMA_signal_1737), .B1_f (new_AGEMA_signal_1738), .Z0_t (stateFF_MUX_inputPar_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_2802), .Z1_t (new_AGEMA_signal_2803), .Z1_f (new_AGEMA_signal_2804) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_27_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_2802), .A1_t (new_AGEMA_signal_2803), .A1_f (new_AGEMA_signal_2804), .B0_t (data_out_s0_t[45]), .B0_f (data_out_s0_f[45]), .B1_t (data_out_s1_t[45]), .B1_f (data_out_s1_f[45]), .Z0_t (stateFF_inputPar[27]), .Z0_f (new_AGEMA_signal_3262), .Z1_t (new_AGEMA_signal_3263), .Z1_f (new_AGEMA_signal_3264) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_XOR1_U1 ( .A0_t (data_out_s0_t[49]), .A0_f (data_out_s0_f[49]), .A1_t (data_out_s1_t[49]), .A1_f (data_out_s1_f[49]), .B0_t (data_in_s0_t[28]), .B0_f (data_in_s0_f[28]), .B1_t (data_in_s1_t[28]), .B1_f (data_in_s1_f[28]), .Z0_t (stateFF_MUX_inputPar_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_1745), .Z1_t (new_AGEMA_signal_1746), .Z1_f (new_AGEMA_signal_1747) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_1745), .B1_t (new_AGEMA_signal_1746), .B1_f (new_AGEMA_signal_1747), .Z0_t (stateFF_MUX_inputPar_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_2805), .Z1_t (new_AGEMA_signal_2806), .Z1_f (new_AGEMA_signal_2807) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_28_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_2805), .A1_t (new_AGEMA_signal_2806), .A1_f (new_AGEMA_signal_2807), .B0_t (data_out_s0_t[49]), .B0_f (data_out_s0_f[49]), .B1_t (data_out_s1_t[49]), .B1_f (data_out_s1_f[49]), .Z0_t (stateFF_inputPar[28]), .Z0_f (new_AGEMA_signal_3265), .Z1_t (new_AGEMA_signal_3266), .Z1_f (new_AGEMA_signal_3267) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_XOR1_U1 ( .A0_t (data_out_s0_t[53]), .A0_f (data_out_s0_f[53]), .A1_t (data_out_s1_t[53]), .A1_f (data_out_s1_f[53]), .B0_t (data_in_s0_t[29]), .B0_f (data_in_s0_f[29]), .B1_t (data_in_s1_t[29]), .B1_f (data_in_s1_f[29]), .Z0_t (stateFF_MUX_inputPar_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_1754), .Z1_t (new_AGEMA_signal_1755), .Z1_f (new_AGEMA_signal_1756) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_1754), .B1_t (new_AGEMA_signal_1755), .B1_f (new_AGEMA_signal_1756), .Z0_t (stateFF_MUX_inputPar_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_2808), .Z1_t (new_AGEMA_signal_2809), .Z1_f (new_AGEMA_signal_2810) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_29_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_2808), .A1_t (new_AGEMA_signal_2809), .A1_f (new_AGEMA_signal_2810), .B0_t (data_out_s0_t[53]), .B0_f (data_out_s0_f[53]), .B1_t (data_out_s1_t[53]), .B1_f (data_out_s1_f[53]), .Z0_t (stateFF_inputPar[29]), .Z0_f (new_AGEMA_signal_3268), .Z1_t (new_AGEMA_signal_3269), .Z1_f (new_AGEMA_signal_3270) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_XOR1_U1 ( .A0_t (data_out_s0_t[57]), .A0_f (data_out_s0_f[57]), .A1_t (data_out_s1_t[57]), .A1_f (data_out_s1_f[57]), .B0_t (data_in_s0_t[30]), .B0_f (data_in_s0_f[30]), .B1_t (data_in_s1_t[30]), .B1_f (data_in_s1_f[30]), .Z0_t (stateFF_MUX_inputPar_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_1763), .Z1_t (new_AGEMA_signal_1764), .Z1_f (new_AGEMA_signal_1765) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_1763), .B1_t (new_AGEMA_signal_1764), .B1_f (new_AGEMA_signal_1765), .Z0_t (stateFF_MUX_inputPar_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_2811), .Z1_t (new_AGEMA_signal_2812), .Z1_f (new_AGEMA_signal_2813) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_30_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_2811), .A1_t (new_AGEMA_signal_2812), .A1_f (new_AGEMA_signal_2813), .B0_t (data_out_s0_t[57]), .B0_f (data_out_s0_f[57]), .B1_t (data_out_s1_t[57]), .B1_f (data_out_s1_f[57]), .Z0_t (stateFF_inputPar[30]), .Z0_f (new_AGEMA_signal_3271), .Z1_t (new_AGEMA_signal_3272), .Z1_f (new_AGEMA_signal_3273) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_XOR1_U1 ( .A0_t (data_out_s0_t[61]), .A0_f (data_out_s0_f[61]), .A1_t (data_out_s1_t[61]), .A1_f (data_out_s1_f[61]), .B0_t (data_in_s0_t[31]), .B0_f (data_in_s0_f[31]), .B1_t (data_in_s1_t[31]), .B1_f (data_in_s1_f[31]), .Z0_t (stateFF_MUX_inputPar_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_1769), .Z1_t (new_AGEMA_signal_1770), .Z1_f (new_AGEMA_signal_1771) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_1769), .B1_t (new_AGEMA_signal_1770), .B1_f (new_AGEMA_signal_1771), .Z0_t (stateFF_MUX_inputPar_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_2814), .Z1_t (new_AGEMA_signal_2815), .Z1_f (new_AGEMA_signal_2816) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_31_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_2814), .A1_t (new_AGEMA_signal_2815), .A1_f (new_AGEMA_signal_2816), .B0_t (data_out_s0_t[61]), .B0_f (data_out_s0_f[61]), .B1_t (data_out_s1_t[61]), .B1_f (data_out_s1_f[61]), .Z0_t (stateFF_inputPar[31]), .Z0_f (new_AGEMA_signal_3274), .Z1_t (new_AGEMA_signal_3275), .Z1_f (new_AGEMA_signal_3276) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_XOR1_U1 ( .A0_t (data_out_s0_t[2]), .A0_f (data_out_s0_f[2]), .A1_t (data_out_s1_t[2]), .A1_f (data_out_s1_f[2]), .B0_t (data_in_s0_t[32]), .B0_f (data_in_s0_f[32]), .B1_t (data_in_s1_t[32]), .B1_f (data_in_s1_f[32]), .Z0_t (stateFF_MUX_inputPar_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_1778), .Z1_t (new_AGEMA_signal_1779), .Z1_f (new_AGEMA_signal_1780) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_1778), .B1_t (new_AGEMA_signal_1779), .B1_f (new_AGEMA_signal_1780), .Z0_t (stateFF_MUX_inputPar_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_2817), .Z1_t (new_AGEMA_signal_2818), .Z1_f (new_AGEMA_signal_2819) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_32_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_2817), .A1_t (new_AGEMA_signal_2818), .A1_f (new_AGEMA_signal_2819), .B0_t (data_out_s0_t[2]), .B0_f (data_out_s0_f[2]), .B1_t (data_out_s1_t[2]), .B1_f (data_out_s1_f[2]), .Z0_t (stateFF_inputPar[32]), .Z0_f (new_AGEMA_signal_3277), .Z1_t (new_AGEMA_signal_3278), .Z1_f (new_AGEMA_signal_3279) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_XOR1_U1 ( .A0_t (data_out_s0_t[6]), .A0_f (data_out_s0_f[6]), .A1_t (data_out_s1_t[6]), .A1_f (data_out_s1_f[6]), .B0_t (data_in_s0_t[33]), .B0_f (data_in_s0_f[33]), .B1_t (data_in_s1_t[33]), .B1_f (data_in_s1_f[33]), .Z0_t (stateFF_MUX_inputPar_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_1787), .Z1_t (new_AGEMA_signal_1788), .Z1_f (new_AGEMA_signal_1789) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_1787), .B1_t (new_AGEMA_signal_1788), .B1_f (new_AGEMA_signal_1789), .Z0_t (stateFF_MUX_inputPar_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_2820), .Z1_t (new_AGEMA_signal_2821), .Z1_f (new_AGEMA_signal_2822) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_33_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_2820), .A1_t (new_AGEMA_signal_2821), .A1_f (new_AGEMA_signal_2822), .B0_t (data_out_s0_t[6]), .B0_f (data_out_s0_f[6]), .B1_t (data_out_s1_t[6]), .B1_f (data_out_s1_f[6]), .Z0_t (stateFF_inputPar[33]), .Z0_f (new_AGEMA_signal_3280), .Z1_t (new_AGEMA_signal_3281), .Z1_f (new_AGEMA_signal_3282) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_XOR1_U1 ( .A0_t (data_out_s0_t[10]), .A0_f (data_out_s0_f[10]), .A1_t (data_out_s1_t[10]), .A1_f (data_out_s1_f[10]), .B0_t (data_in_s0_t[34]), .B0_f (data_in_s0_f[34]), .B1_t (data_in_s1_t[34]), .B1_f (data_in_s1_f[34]), .Z0_t (stateFF_MUX_inputPar_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_1796), .Z1_t (new_AGEMA_signal_1797), .Z1_f (new_AGEMA_signal_1798) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_1796), .B1_t (new_AGEMA_signal_1797), .B1_f (new_AGEMA_signal_1798), .Z0_t (stateFF_MUX_inputPar_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_2823), .Z1_t (new_AGEMA_signal_2824), .Z1_f (new_AGEMA_signal_2825) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_34_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_2823), .A1_t (new_AGEMA_signal_2824), .A1_f (new_AGEMA_signal_2825), .B0_t (data_out_s0_t[10]), .B0_f (data_out_s0_f[10]), .B1_t (data_out_s1_t[10]), .B1_f (data_out_s1_f[10]), .Z0_t (stateFF_inputPar[34]), .Z0_f (new_AGEMA_signal_3283), .Z1_t (new_AGEMA_signal_3284), .Z1_f (new_AGEMA_signal_3285) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_XOR1_U1 ( .A0_t (data_out_s0_t[14]), .A0_f (data_out_s0_f[14]), .A1_t (data_out_s1_t[14]), .A1_f (data_out_s1_f[14]), .B0_t (data_in_s0_t[35]), .B0_f (data_in_s0_f[35]), .B1_t (data_in_s1_t[35]), .B1_f (data_in_s1_f[35]), .Z0_t (stateFF_MUX_inputPar_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_1805), .Z1_t (new_AGEMA_signal_1806), .Z1_f (new_AGEMA_signal_1807) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_1805), .B1_t (new_AGEMA_signal_1806), .B1_f (new_AGEMA_signal_1807), .Z0_t (stateFF_MUX_inputPar_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_2826), .Z1_t (new_AGEMA_signal_2827), .Z1_f (new_AGEMA_signal_2828) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_35_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_2826), .A1_t (new_AGEMA_signal_2827), .A1_f (new_AGEMA_signal_2828), .B0_t (data_out_s0_t[14]), .B0_f (data_out_s0_f[14]), .B1_t (data_out_s1_t[14]), .B1_f (data_out_s1_f[14]), .Z0_t (stateFF_inputPar[35]), .Z0_f (new_AGEMA_signal_3286), .Z1_t (new_AGEMA_signal_3287), .Z1_f (new_AGEMA_signal_3288) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_XOR1_U1 ( .A0_t (data_out_s0_t[18]), .A0_f (data_out_s0_f[18]), .A1_t (data_out_s1_t[18]), .A1_f (data_out_s1_f[18]), .B0_t (data_in_s0_t[36]), .B0_f (data_in_s0_f[36]), .B1_t (data_in_s1_t[36]), .B1_f (data_in_s1_f[36]), .Z0_t (stateFF_MUX_inputPar_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_1814), .Z1_t (new_AGEMA_signal_1815), .Z1_f (new_AGEMA_signal_1816) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_1814), .B1_t (new_AGEMA_signal_1815), .B1_f (new_AGEMA_signal_1816), .Z0_t (stateFF_MUX_inputPar_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_2829), .Z1_t (new_AGEMA_signal_2830), .Z1_f (new_AGEMA_signal_2831) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_36_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_2829), .A1_t (new_AGEMA_signal_2830), .A1_f (new_AGEMA_signal_2831), .B0_t (data_out_s0_t[18]), .B0_f (data_out_s0_f[18]), .B1_t (data_out_s1_t[18]), .B1_f (data_out_s1_f[18]), .Z0_t (stateFF_inputPar[36]), .Z0_f (new_AGEMA_signal_3289), .Z1_t (new_AGEMA_signal_3290), .Z1_f (new_AGEMA_signal_3291) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_XOR1_U1 ( .A0_t (data_out_s0_t[22]), .A0_f (data_out_s0_f[22]), .A1_t (data_out_s1_t[22]), .A1_f (data_out_s1_f[22]), .B0_t (data_in_s0_t[37]), .B0_f (data_in_s0_f[37]), .B1_t (data_in_s1_t[37]), .B1_f (data_in_s1_f[37]), .Z0_t (stateFF_MUX_inputPar_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_1823), .Z1_t (new_AGEMA_signal_1824), .Z1_f (new_AGEMA_signal_1825) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_1823), .B1_t (new_AGEMA_signal_1824), .B1_f (new_AGEMA_signal_1825), .Z0_t (stateFF_MUX_inputPar_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_2832), .Z1_t (new_AGEMA_signal_2833), .Z1_f (new_AGEMA_signal_2834) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_37_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_2832), .A1_t (new_AGEMA_signal_2833), .A1_f (new_AGEMA_signal_2834), .B0_t (data_out_s0_t[22]), .B0_f (data_out_s0_f[22]), .B1_t (data_out_s1_t[22]), .B1_f (data_out_s1_f[22]), .Z0_t (stateFF_inputPar[37]), .Z0_f (new_AGEMA_signal_3292), .Z1_t (new_AGEMA_signal_3293), .Z1_f (new_AGEMA_signal_3294) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_XOR1_U1 ( .A0_t (data_out_s0_t[26]), .A0_f (data_out_s0_f[26]), .A1_t (data_out_s1_t[26]), .A1_f (data_out_s1_f[26]), .B0_t (data_in_s0_t[38]), .B0_f (data_in_s0_f[38]), .B1_t (data_in_s1_t[38]), .B1_f (data_in_s1_f[38]), .Z0_t (stateFF_MUX_inputPar_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_1832), .Z1_t (new_AGEMA_signal_1833), .Z1_f (new_AGEMA_signal_1834) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_1832), .B1_t (new_AGEMA_signal_1833), .B1_f (new_AGEMA_signal_1834), .Z0_t (stateFF_MUX_inputPar_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_2835), .Z1_t (new_AGEMA_signal_2836), .Z1_f (new_AGEMA_signal_2837) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_38_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_2835), .A1_t (new_AGEMA_signal_2836), .A1_f (new_AGEMA_signal_2837), .B0_t (data_out_s0_t[26]), .B0_f (data_out_s0_f[26]), .B1_t (data_out_s1_t[26]), .B1_f (data_out_s1_f[26]), .Z0_t (stateFF_inputPar[38]), .Z0_f (new_AGEMA_signal_3295), .Z1_t (new_AGEMA_signal_3296), .Z1_f (new_AGEMA_signal_3297) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_XOR1_U1 ( .A0_t (data_out_s0_t[30]), .A0_f (data_out_s0_f[30]), .A1_t (data_out_s1_t[30]), .A1_f (data_out_s1_f[30]), .B0_t (data_in_s0_t[39]), .B0_f (data_in_s0_f[39]), .B1_t (data_in_s1_t[39]), .B1_f (data_in_s1_f[39]), .Z0_t (stateFF_MUX_inputPar_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_1841), .Z1_t (new_AGEMA_signal_1842), .Z1_f (new_AGEMA_signal_1843) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_1841), .B1_t (new_AGEMA_signal_1842), .B1_f (new_AGEMA_signal_1843), .Z0_t (stateFF_MUX_inputPar_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_2838), .Z1_t (new_AGEMA_signal_2839), .Z1_f (new_AGEMA_signal_2840) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_39_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_2838), .A1_t (new_AGEMA_signal_2839), .A1_f (new_AGEMA_signal_2840), .B0_t (data_out_s0_t[30]), .B0_f (data_out_s0_f[30]), .B1_t (data_out_s1_t[30]), .B1_f (data_out_s1_f[30]), .Z0_t (stateFF_inputPar[39]), .Z0_f (new_AGEMA_signal_3298), .Z1_t (new_AGEMA_signal_3299), .Z1_f (new_AGEMA_signal_3300) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_XOR1_U1 ( .A0_t (data_out_s0_t[34]), .A0_f (data_out_s0_f[34]), .A1_t (data_out_s1_t[34]), .A1_f (data_out_s1_f[34]), .B0_t (data_in_s0_t[40]), .B0_f (data_in_s0_f[40]), .B1_t (data_in_s1_t[40]), .B1_f (data_in_s1_f[40]), .Z0_t (stateFF_MUX_inputPar_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_1850), .Z1_t (new_AGEMA_signal_1851), .Z1_f (new_AGEMA_signal_1852) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_1850), .B1_t (new_AGEMA_signal_1851), .B1_f (new_AGEMA_signal_1852), .Z0_t (stateFF_MUX_inputPar_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_2841), .Z1_t (new_AGEMA_signal_2842), .Z1_f (new_AGEMA_signal_2843) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_40_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_2841), .A1_t (new_AGEMA_signal_2842), .A1_f (new_AGEMA_signal_2843), .B0_t (data_out_s0_t[34]), .B0_f (data_out_s0_f[34]), .B1_t (data_out_s1_t[34]), .B1_f (data_out_s1_f[34]), .Z0_t (stateFF_inputPar[40]), .Z0_f (new_AGEMA_signal_3301), .Z1_t (new_AGEMA_signal_3302), .Z1_f (new_AGEMA_signal_3303) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_XOR1_U1 ( .A0_t (data_out_s0_t[38]), .A0_f (data_out_s0_f[38]), .A1_t (data_out_s1_t[38]), .A1_f (data_out_s1_f[38]), .B0_t (data_in_s0_t[41]), .B0_f (data_in_s0_f[41]), .B1_t (data_in_s1_t[41]), .B1_f (data_in_s1_f[41]), .Z0_t (stateFF_MUX_inputPar_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_1859), .Z1_t (new_AGEMA_signal_1860), .Z1_f (new_AGEMA_signal_1861) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_1859), .B1_t (new_AGEMA_signal_1860), .B1_f (new_AGEMA_signal_1861), .Z0_t (stateFF_MUX_inputPar_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_2844), .Z1_t (new_AGEMA_signal_2845), .Z1_f (new_AGEMA_signal_2846) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_41_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_2844), .A1_t (new_AGEMA_signal_2845), .A1_f (new_AGEMA_signal_2846), .B0_t (data_out_s0_t[38]), .B0_f (data_out_s0_f[38]), .B1_t (data_out_s1_t[38]), .B1_f (data_out_s1_f[38]), .Z0_t (stateFF_inputPar[41]), .Z0_f (new_AGEMA_signal_3304), .Z1_t (new_AGEMA_signal_3305), .Z1_f (new_AGEMA_signal_3306) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_XOR1_U1 ( .A0_t (data_out_s0_t[42]), .A0_f (data_out_s0_f[42]), .A1_t (data_out_s1_t[42]), .A1_f (data_out_s1_f[42]), .B0_t (data_in_s0_t[42]), .B0_f (data_in_s0_f[42]), .B1_t (data_in_s1_t[42]), .B1_f (data_in_s1_f[42]), .Z0_t (stateFF_MUX_inputPar_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_1868), .Z1_t (new_AGEMA_signal_1869), .Z1_f (new_AGEMA_signal_1870) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_1868), .B1_t (new_AGEMA_signal_1869), .B1_f (new_AGEMA_signal_1870), .Z0_t (stateFF_MUX_inputPar_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_2847), .Z1_t (new_AGEMA_signal_2848), .Z1_f (new_AGEMA_signal_2849) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_42_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_2847), .A1_t (new_AGEMA_signal_2848), .A1_f (new_AGEMA_signal_2849), .B0_t (data_out_s0_t[42]), .B0_f (data_out_s0_f[42]), .B1_t (data_out_s1_t[42]), .B1_f (data_out_s1_f[42]), .Z0_t (stateFF_inputPar[42]), .Z0_f (new_AGEMA_signal_3307), .Z1_t (new_AGEMA_signal_3308), .Z1_f (new_AGEMA_signal_3309) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_XOR1_U1 ( .A0_t (data_out_s0_t[46]), .A0_f (data_out_s0_f[46]), .A1_t (data_out_s1_t[46]), .A1_f (data_out_s1_f[46]), .B0_t (data_in_s0_t[43]), .B0_f (data_in_s0_f[43]), .B1_t (data_in_s1_t[43]), .B1_f (data_in_s1_f[43]), .Z0_t (stateFF_MUX_inputPar_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_1877), .Z1_t (new_AGEMA_signal_1878), .Z1_f (new_AGEMA_signal_1879) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_1877), .B1_t (new_AGEMA_signal_1878), .B1_f (new_AGEMA_signal_1879), .Z0_t (stateFF_MUX_inputPar_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_2850), .Z1_t (new_AGEMA_signal_2851), .Z1_f (new_AGEMA_signal_2852) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_43_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_2850), .A1_t (new_AGEMA_signal_2851), .A1_f (new_AGEMA_signal_2852), .B0_t (data_out_s0_t[46]), .B0_f (data_out_s0_f[46]), .B1_t (data_out_s1_t[46]), .B1_f (data_out_s1_f[46]), .Z0_t (stateFF_inputPar[43]), .Z0_f (new_AGEMA_signal_3310), .Z1_t (new_AGEMA_signal_3311), .Z1_f (new_AGEMA_signal_3312) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_XOR1_U1 ( .A0_t (data_out_s0_t[50]), .A0_f (data_out_s0_f[50]), .A1_t (data_out_s1_t[50]), .A1_f (data_out_s1_f[50]), .B0_t (data_in_s0_t[44]), .B0_f (data_in_s0_f[44]), .B1_t (data_in_s1_t[44]), .B1_f (data_in_s1_f[44]), .Z0_t (stateFF_MUX_inputPar_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_1886), .Z1_t (new_AGEMA_signal_1887), .Z1_f (new_AGEMA_signal_1888) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_1886), .B1_t (new_AGEMA_signal_1887), .B1_f (new_AGEMA_signal_1888), .Z0_t (stateFF_MUX_inputPar_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_2853), .Z1_t (new_AGEMA_signal_2854), .Z1_f (new_AGEMA_signal_2855) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_44_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_2853), .A1_t (new_AGEMA_signal_2854), .A1_f (new_AGEMA_signal_2855), .B0_t (data_out_s0_t[50]), .B0_f (data_out_s0_f[50]), .B1_t (data_out_s1_t[50]), .B1_f (data_out_s1_f[50]), .Z0_t (stateFF_inputPar[44]), .Z0_f (new_AGEMA_signal_3313), .Z1_t (new_AGEMA_signal_3314), .Z1_f (new_AGEMA_signal_3315) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_XOR1_U1 ( .A0_t (data_out_s0_t[54]), .A0_f (data_out_s0_f[54]), .A1_t (data_out_s1_t[54]), .A1_f (data_out_s1_f[54]), .B0_t (data_in_s0_t[45]), .B0_f (data_in_s0_f[45]), .B1_t (data_in_s1_t[45]), .B1_f (data_in_s1_f[45]), .Z0_t (stateFF_MUX_inputPar_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_1895), .Z1_t (new_AGEMA_signal_1896), .Z1_f (new_AGEMA_signal_1897) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_1895), .B1_t (new_AGEMA_signal_1896), .B1_f (new_AGEMA_signal_1897), .Z0_t (stateFF_MUX_inputPar_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_2856), .Z1_t (new_AGEMA_signal_2857), .Z1_f (new_AGEMA_signal_2858) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_45_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_2856), .A1_t (new_AGEMA_signal_2857), .A1_f (new_AGEMA_signal_2858), .B0_t (data_out_s0_t[54]), .B0_f (data_out_s0_f[54]), .B1_t (data_out_s1_t[54]), .B1_f (data_out_s1_f[54]), .Z0_t (stateFF_inputPar[45]), .Z0_f (new_AGEMA_signal_3316), .Z1_t (new_AGEMA_signal_3317), .Z1_f (new_AGEMA_signal_3318) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_XOR1_U1 ( .A0_t (data_out_s0_t[58]), .A0_f (data_out_s0_f[58]), .A1_t (data_out_s1_t[58]), .A1_f (data_out_s1_f[58]), .B0_t (data_in_s0_t[46]), .B0_f (data_in_s0_f[46]), .B1_t (data_in_s1_t[46]), .B1_f (data_in_s1_f[46]), .Z0_t (stateFF_MUX_inputPar_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_1904), .Z1_t (new_AGEMA_signal_1905), .Z1_f (new_AGEMA_signal_1906) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_1904), .B1_t (new_AGEMA_signal_1905), .B1_f (new_AGEMA_signal_1906), .Z0_t (stateFF_MUX_inputPar_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_2859), .Z1_t (new_AGEMA_signal_2860), .Z1_f (new_AGEMA_signal_2861) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_46_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_2859), .A1_t (new_AGEMA_signal_2860), .A1_f (new_AGEMA_signal_2861), .B0_t (data_out_s0_t[58]), .B0_f (data_out_s0_f[58]), .B1_t (data_out_s1_t[58]), .B1_f (data_out_s1_f[58]), .Z0_t (stateFF_inputPar[46]), .Z0_f (new_AGEMA_signal_3319), .Z1_t (new_AGEMA_signal_3320), .Z1_f (new_AGEMA_signal_3321) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_XOR1_U1 ( .A0_t (data_out_s0_t[62]), .A0_f (data_out_s0_f[62]), .A1_t (data_out_s1_t[62]), .A1_f (data_out_s1_f[62]), .B0_t (data_in_s0_t[47]), .B0_f (data_in_s0_f[47]), .B1_t (data_in_s1_t[47]), .B1_f (data_in_s1_f[47]), .Z0_t (stateFF_MUX_inputPar_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_1910), .Z1_t (new_AGEMA_signal_1911), .Z1_f (new_AGEMA_signal_1912) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_1910), .B1_t (new_AGEMA_signal_1911), .B1_f (new_AGEMA_signal_1912), .Z0_t (stateFF_MUX_inputPar_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_2862), .Z1_t (new_AGEMA_signal_2863), .Z1_f (new_AGEMA_signal_2864) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_47_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_2862), .A1_t (new_AGEMA_signal_2863), .A1_f (new_AGEMA_signal_2864), .B0_t (data_out_s0_t[62]), .B0_f (data_out_s0_f[62]), .B1_t (data_out_s1_t[62]), .B1_f (data_out_s1_f[62]), .Z0_t (stateFF_inputPar[47]), .Z0_f (new_AGEMA_signal_3322), .Z1_t (new_AGEMA_signal_3323), .Z1_f (new_AGEMA_signal_3324) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_XOR1_U1 ( .A0_t (data_out_s0_t[3]), .A0_f (data_out_s0_f[3]), .A1_t (data_out_s1_t[3]), .A1_f (data_out_s1_f[3]), .B0_t (data_in_s0_t[48]), .B0_f (data_in_s0_f[48]), .B1_t (data_in_s1_t[48]), .B1_f (data_in_s1_f[48]), .Z0_t (stateFF_MUX_inputPar_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_1919), .Z1_t (new_AGEMA_signal_1920), .Z1_f (new_AGEMA_signal_1921) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_1919), .B1_t (new_AGEMA_signal_1920), .B1_f (new_AGEMA_signal_1921), .Z0_t (stateFF_MUX_inputPar_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_2865), .Z1_t (new_AGEMA_signal_2866), .Z1_f (new_AGEMA_signal_2867) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_48_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_2865), .A1_t (new_AGEMA_signal_2866), .A1_f (new_AGEMA_signal_2867), .B0_t (data_out_s0_t[3]), .B0_f (data_out_s0_f[3]), .B1_t (data_out_s1_t[3]), .B1_f (data_out_s1_f[3]), .Z0_t (stateFF_inputPar[48]), .Z0_f (new_AGEMA_signal_3325), .Z1_t (new_AGEMA_signal_3326), .Z1_f (new_AGEMA_signal_3327) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_XOR1_U1 ( .A0_t (data_out_s0_t[7]), .A0_f (data_out_s0_f[7]), .A1_t (data_out_s1_t[7]), .A1_f (data_out_s1_f[7]), .B0_t (data_in_s0_t[49]), .B0_f (data_in_s0_f[49]), .B1_t (data_in_s1_t[49]), .B1_f (data_in_s1_f[49]), .Z0_t (stateFF_MUX_inputPar_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_1928), .Z1_t (new_AGEMA_signal_1929), .Z1_f (new_AGEMA_signal_1930) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_1928), .B1_t (new_AGEMA_signal_1929), .B1_f (new_AGEMA_signal_1930), .Z0_t (stateFF_MUX_inputPar_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_2868), .Z1_t (new_AGEMA_signal_2869), .Z1_f (new_AGEMA_signal_2870) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_49_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_2868), .A1_t (new_AGEMA_signal_2869), .A1_f (new_AGEMA_signal_2870), .B0_t (data_out_s0_t[7]), .B0_f (data_out_s0_f[7]), .B1_t (data_out_s1_t[7]), .B1_f (data_out_s1_f[7]), .Z0_t (stateFF_inputPar[49]), .Z0_f (new_AGEMA_signal_3328), .Z1_t (new_AGEMA_signal_3329), .Z1_f (new_AGEMA_signal_3330) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_XOR1_U1 ( .A0_t (data_out_s0_t[11]), .A0_f (data_out_s0_f[11]), .A1_t (data_out_s1_t[11]), .A1_f (data_out_s1_f[11]), .B0_t (data_in_s0_t[50]), .B0_f (data_in_s0_f[50]), .B1_t (data_in_s1_t[50]), .B1_f (data_in_s1_f[50]), .Z0_t (stateFF_MUX_inputPar_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_1937), .Z1_t (new_AGEMA_signal_1938), .Z1_f (new_AGEMA_signal_1939) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_1937), .B1_t (new_AGEMA_signal_1938), .B1_f (new_AGEMA_signal_1939), .Z0_t (stateFF_MUX_inputPar_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_2871), .Z1_t (new_AGEMA_signal_2872), .Z1_f (new_AGEMA_signal_2873) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_50_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_2871), .A1_t (new_AGEMA_signal_2872), .A1_f (new_AGEMA_signal_2873), .B0_t (data_out_s0_t[11]), .B0_f (data_out_s0_f[11]), .B1_t (data_out_s1_t[11]), .B1_f (data_out_s1_f[11]), .Z0_t (stateFF_inputPar[50]), .Z0_f (new_AGEMA_signal_3331), .Z1_t (new_AGEMA_signal_3332), .Z1_f (new_AGEMA_signal_3333) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_XOR1_U1 ( .A0_t (data_out_s0_t[15]), .A0_f (data_out_s0_f[15]), .A1_t (data_out_s1_t[15]), .A1_f (data_out_s1_f[15]), .B0_t (data_in_s0_t[51]), .B0_f (data_in_s0_f[51]), .B1_t (data_in_s1_t[51]), .B1_f (data_in_s1_f[51]), .Z0_t (stateFF_MUX_inputPar_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_1946), .Z1_t (new_AGEMA_signal_1947), .Z1_f (new_AGEMA_signal_1948) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_1946), .B1_t (new_AGEMA_signal_1947), .B1_f (new_AGEMA_signal_1948), .Z0_t (stateFF_MUX_inputPar_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_2874), .Z1_t (new_AGEMA_signal_2875), .Z1_f (new_AGEMA_signal_2876) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_51_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_2874), .A1_t (new_AGEMA_signal_2875), .A1_f (new_AGEMA_signal_2876), .B0_t (data_out_s0_t[15]), .B0_f (data_out_s0_f[15]), .B1_t (data_out_s1_t[15]), .B1_f (data_out_s1_f[15]), .Z0_t (stateFF_inputPar[51]), .Z0_f (new_AGEMA_signal_3334), .Z1_t (new_AGEMA_signal_3335), .Z1_f (new_AGEMA_signal_3336) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_XOR1_U1 ( .A0_t (data_out_s0_t[19]), .A0_f (data_out_s0_f[19]), .A1_t (data_out_s1_t[19]), .A1_f (data_out_s1_f[19]), .B0_t (data_in_s0_t[52]), .B0_f (data_in_s0_f[52]), .B1_t (data_in_s1_t[52]), .B1_f (data_in_s1_f[52]), .Z0_t (stateFF_MUX_inputPar_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_1955), .Z1_t (new_AGEMA_signal_1956), .Z1_f (new_AGEMA_signal_1957) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_1955), .B1_t (new_AGEMA_signal_1956), .B1_f (new_AGEMA_signal_1957), .Z0_t (stateFF_MUX_inputPar_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_2877), .Z1_t (new_AGEMA_signal_2878), .Z1_f (new_AGEMA_signal_2879) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_52_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_2877), .A1_t (new_AGEMA_signal_2878), .A1_f (new_AGEMA_signal_2879), .B0_t (data_out_s0_t[19]), .B0_f (data_out_s0_f[19]), .B1_t (data_out_s1_t[19]), .B1_f (data_out_s1_f[19]), .Z0_t (stateFF_inputPar[52]), .Z0_f (new_AGEMA_signal_3337), .Z1_t (new_AGEMA_signal_3338), .Z1_f (new_AGEMA_signal_3339) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_XOR1_U1 ( .A0_t (data_out_s0_t[23]), .A0_f (data_out_s0_f[23]), .A1_t (data_out_s1_t[23]), .A1_f (data_out_s1_f[23]), .B0_t (data_in_s0_t[53]), .B0_f (data_in_s0_f[53]), .B1_t (data_in_s1_t[53]), .B1_f (data_in_s1_f[53]), .Z0_t (stateFF_MUX_inputPar_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_1964), .Z1_t (new_AGEMA_signal_1965), .Z1_f (new_AGEMA_signal_1966) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_1964), .B1_t (new_AGEMA_signal_1965), .B1_f (new_AGEMA_signal_1966), .Z0_t (stateFF_MUX_inputPar_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_2880), .Z1_t (new_AGEMA_signal_2881), .Z1_f (new_AGEMA_signal_2882) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_53_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_2880), .A1_t (new_AGEMA_signal_2881), .A1_f (new_AGEMA_signal_2882), .B0_t (data_out_s0_t[23]), .B0_f (data_out_s0_f[23]), .B1_t (data_out_s1_t[23]), .B1_f (data_out_s1_f[23]), .Z0_t (stateFF_inputPar[53]), .Z0_f (new_AGEMA_signal_3340), .Z1_t (new_AGEMA_signal_3341), .Z1_f (new_AGEMA_signal_3342) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_XOR1_U1 ( .A0_t (data_out_s0_t[27]), .A0_f (data_out_s0_f[27]), .A1_t (data_out_s1_t[27]), .A1_f (data_out_s1_f[27]), .B0_t (data_in_s0_t[54]), .B0_f (data_in_s0_f[54]), .B1_t (data_in_s1_t[54]), .B1_f (data_in_s1_f[54]), .Z0_t (stateFF_MUX_inputPar_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_1973), .Z1_t (new_AGEMA_signal_1974), .Z1_f (new_AGEMA_signal_1975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_1973), .B1_t (new_AGEMA_signal_1974), .B1_f (new_AGEMA_signal_1975), .Z0_t (stateFF_MUX_inputPar_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_2883), .Z1_t (new_AGEMA_signal_2884), .Z1_f (new_AGEMA_signal_2885) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_54_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_2883), .A1_t (new_AGEMA_signal_2884), .A1_f (new_AGEMA_signal_2885), .B0_t (data_out_s0_t[27]), .B0_f (data_out_s0_f[27]), .B1_t (data_out_s1_t[27]), .B1_f (data_out_s1_f[27]), .Z0_t (stateFF_inputPar[54]), .Z0_f (new_AGEMA_signal_3343), .Z1_t (new_AGEMA_signal_3344), .Z1_f (new_AGEMA_signal_3345) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_XOR1_U1 ( .A0_t (data_out_s0_t[31]), .A0_f (data_out_s0_f[31]), .A1_t (data_out_s1_t[31]), .A1_f (data_out_s1_f[31]), .B0_t (data_in_s0_t[55]), .B0_f (data_in_s0_f[55]), .B1_t (data_in_s1_t[55]), .B1_f (data_in_s1_f[55]), .Z0_t (stateFF_MUX_inputPar_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_1982), .Z1_t (new_AGEMA_signal_1983), .Z1_f (new_AGEMA_signal_1984) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_1982), .B1_t (new_AGEMA_signal_1983), .B1_f (new_AGEMA_signal_1984), .Z0_t (stateFF_MUX_inputPar_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_2886), .Z1_t (new_AGEMA_signal_2887), .Z1_f (new_AGEMA_signal_2888) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_55_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_2886), .A1_t (new_AGEMA_signal_2887), .A1_f (new_AGEMA_signal_2888), .B0_t (data_out_s0_t[31]), .B0_f (data_out_s0_f[31]), .B1_t (data_out_s1_t[31]), .B1_f (data_out_s1_f[31]), .Z0_t (stateFF_inputPar[55]), .Z0_f (new_AGEMA_signal_3346), .Z1_t (new_AGEMA_signal_3347), .Z1_f (new_AGEMA_signal_3348) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_XOR1_U1 ( .A0_t (data_out_s0_t[35]), .A0_f (data_out_s0_f[35]), .A1_t (data_out_s1_t[35]), .A1_f (data_out_s1_f[35]), .B0_t (data_in_s0_t[56]), .B0_f (data_in_s0_f[56]), .B1_t (data_in_s1_t[56]), .B1_f (data_in_s1_f[56]), .Z0_t (stateFF_MUX_inputPar_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_1991), .Z1_t (new_AGEMA_signal_1992), .Z1_f (new_AGEMA_signal_1993) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_1991), .B1_t (new_AGEMA_signal_1992), .B1_f (new_AGEMA_signal_1993), .Z0_t (stateFF_MUX_inputPar_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_2889), .Z1_t (new_AGEMA_signal_2890), .Z1_f (new_AGEMA_signal_2891) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_56_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_2889), .A1_t (new_AGEMA_signal_2890), .A1_f (new_AGEMA_signal_2891), .B0_t (data_out_s0_t[35]), .B0_f (data_out_s0_f[35]), .B1_t (data_out_s1_t[35]), .B1_f (data_out_s1_f[35]), .Z0_t (stateFF_inputPar[56]), .Z0_f (new_AGEMA_signal_3349), .Z1_t (new_AGEMA_signal_3350), .Z1_f (new_AGEMA_signal_3351) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_XOR1_U1 ( .A0_t (data_out_s0_t[39]), .A0_f (data_out_s0_f[39]), .A1_t (data_out_s1_t[39]), .A1_f (data_out_s1_f[39]), .B0_t (data_in_s0_t[57]), .B0_f (data_in_s0_f[57]), .B1_t (data_in_s1_t[57]), .B1_f (data_in_s1_f[57]), .Z0_t (stateFF_MUX_inputPar_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_2000), .Z1_t (new_AGEMA_signal_2001), .Z1_f (new_AGEMA_signal_2002) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_2000), .B1_t (new_AGEMA_signal_2001), .B1_f (new_AGEMA_signal_2002), .Z0_t (stateFF_MUX_inputPar_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_2892), .Z1_t (new_AGEMA_signal_2893), .Z1_f (new_AGEMA_signal_2894) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_57_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_2892), .A1_t (new_AGEMA_signal_2893), .A1_f (new_AGEMA_signal_2894), .B0_t (data_out_s0_t[39]), .B0_f (data_out_s0_f[39]), .B1_t (data_out_s1_t[39]), .B1_f (data_out_s1_f[39]), .Z0_t (stateFF_inputPar[57]), .Z0_f (new_AGEMA_signal_3352), .Z1_t (new_AGEMA_signal_3353), .Z1_f (new_AGEMA_signal_3354) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_XOR1_U1 ( .A0_t (data_out_s0_t[43]), .A0_f (data_out_s0_f[43]), .A1_t (data_out_s1_t[43]), .A1_f (data_out_s1_f[43]), .B0_t (data_in_s0_t[58]), .B0_f (data_in_s0_f[58]), .B1_t (data_in_s1_t[58]), .B1_f (data_in_s1_f[58]), .Z0_t (stateFF_MUX_inputPar_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_2009), .Z1_t (new_AGEMA_signal_2010), .Z1_f (new_AGEMA_signal_2011) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_2009), .B1_t (new_AGEMA_signal_2010), .B1_f (new_AGEMA_signal_2011), .Z0_t (stateFF_MUX_inputPar_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_2895), .Z1_t (new_AGEMA_signal_2896), .Z1_f (new_AGEMA_signal_2897) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_58_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_2895), .A1_t (new_AGEMA_signal_2896), .A1_f (new_AGEMA_signal_2897), .B0_t (data_out_s0_t[43]), .B0_f (data_out_s0_f[43]), .B1_t (data_out_s1_t[43]), .B1_f (data_out_s1_f[43]), .Z0_t (stateFF_inputPar[58]), .Z0_f (new_AGEMA_signal_3355), .Z1_t (new_AGEMA_signal_3356), .Z1_f (new_AGEMA_signal_3357) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_XOR1_U1 ( .A0_t (data_out_s0_t[47]), .A0_f (data_out_s0_f[47]), .A1_t (data_out_s1_t[47]), .A1_f (data_out_s1_f[47]), .B0_t (data_in_s0_t[59]), .B0_f (data_in_s0_f[59]), .B1_t (data_in_s1_t[59]), .B1_f (data_in_s1_f[59]), .Z0_t (stateFF_MUX_inputPar_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_2018), .Z1_t (new_AGEMA_signal_2019), .Z1_f (new_AGEMA_signal_2020) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_2018), .B1_t (new_AGEMA_signal_2019), .B1_f (new_AGEMA_signal_2020), .Z0_t (stateFF_MUX_inputPar_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_2898), .Z1_t (new_AGEMA_signal_2899), .Z1_f (new_AGEMA_signal_2900) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_59_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_2898), .A1_t (new_AGEMA_signal_2899), .A1_f (new_AGEMA_signal_2900), .B0_t (data_out_s0_t[47]), .B0_f (data_out_s0_f[47]), .B1_t (data_out_s1_t[47]), .B1_f (data_out_s1_f[47]), .Z0_t (stateFF_inputPar[59]), .Z0_f (new_AGEMA_signal_3358), .Z1_t (new_AGEMA_signal_3359), .Z1_f (new_AGEMA_signal_3360) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_XOR1_U1 ( .A0_t (data_out_s0_t[51]), .A0_f (data_out_s0_f[51]), .A1_t (data_out_s1_t[51]), .A1_f (data_out_s1_f[51]), .B0_t (data_in_s0_t[60]), .B0_f (data_in_s0_f[60]), .B1_t (data_in_s1_t[60]), .B1_f (data_in_s1_f[60]), .Z0_t (stateFF_MUX_inputPar_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_2027), .Z1_t (new_AGEMA_signal_2028), .Z1_f (new_AGEMA_signal_2029) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_2027), .B1_t (new_AGEMA_signal_2028), .B1_f (new_AGEMA_signal_2029), .Z0_t (stateFF_MUX_inputPar_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_2901), .Z1_t (new_AGEMA_signal_2902), .Z1_f (new_AGEMA_signal_2903) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_60_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_2901), .A1_t (new_AGEMA_signal_2902), .A1_f (new_AGEMA_signal_2903), .B0_t (data_out_s0_t[51]), .B0_f (data_out_s0_f[51]), .B1_t (data_out_s1_t[51]), .B1_f (data_out_s1_f[51]), .Z0_t (stateFF_inputPar[60]), .Z0_f (new_AGEMA_signal_3361), .Z1_t (new_AGEMA_signal_3362), .Z1_f (new_AGEMA_signal_3363) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_XOR1_U1 ( .A0_t (data_out_s0_t[55]), .A0_f (data_out_s0_f[55]), .A1_t (data_out_s1_t[55]), .A1_f (data_out_s1_f[55]), .B0_t (data_in_s0_t[61]), .B0_f (data_in_s0_f[61]), .B1_t (data_in_s1_t[61]), .B1_f (data_in_s1_f[61]), .Z0_t (stateFF_MUX_inputPar_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_2036), .Z1_t (new_AGEMA_signal_2037), .Z1_f (new_AGEMA_signal_2038) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_2036), .B1_t (new_AGEMA_signal_2037), .B1_f (new_AGEMA_signal_2038), .Z0_t (stateFF_MUX_inputPar_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_2904), .Z1_t (new_AGEMA_signal_2905), .Z1_f (new_AGEMA_signal_2906) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_61_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_2904), .A1_t (new_AGEMA_signal_2905), .A1_f (new_AGEMA_signal_2906), .B0_t (data_out_s0_t[55]), .B0_f (data_out_s0_f[55]), .B1_t (data_out_s1_t[55]), .B1_f (data_out_s1_f[55]), .Z0_t (stateFF_inputPar[61]), .Z0_f (new_AGEMA_signal_3364), .Z1_t (new_AGEMA_signal_3365), .Z1_f (new_AGEMA_signal_3366) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_XOR1_U1 ( .A0_t (data_out_s0_t[59]), .A0_f (data_out_s0_f[59]), .A1_t (data_out_s1_t[59]), .A1_f (data_out_s1_f[59]), .B0_t (data_in_s0_t[62]), .B0_f (data_in_s0_f[62]), .B1_t (data_in_s1_t[62]), .B1_f (data_in_s1_f[62]), .Z0_t (stateFF_MUX_inputPar_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_2045), .Z1_t (new_AGEMA_signal_2046), .Z1_f (new_AGEMA_signal_2047) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_2045), .B1_t (new_AGEMA_signal_2046), .B1_f (new_AGEMA_signal_2047), .Z0_t (stateFF_MUX_inputPar_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_2907), .Z1_t (new_AGEMA_signal_2908), .Z1_f (new_AGEMA_signal_2909) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_62_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_2907), .A1_t (new_AGEMA_signal_2908), .A1_f (new_AGEMA_signal_2909), .B0_t (data_out_s0_t[59]), .B0_f (data_out_s0_f[59]), .B1_t (data_out_s1_t[59]), .B1_f (data_out_s1_f[59]), .Z0_t (stateFF_inputPar[62]), .Z0_f (new_AGEMA_signal_3367), .Z1_t (new_AGEMA_signal_3368), .Z1_f (new_AGEMA_signal_3369) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_XOR1_U1 ( .A0_t (data_out_s0_t[63]), .A0_f (data_out_s0_f[63]), .A1_t (data_out_s1_t[63]), .A1_f (data_out_s1_f[63]), .B0_t (data_in_s0_t[63]), .B0_f (data_in_s0_f[63]), .B1_t (data_in_s1_t[63]), .B1_f (data_in_s1_f[63]), .Z0_t (stateFF_MUX_inputPar_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_2051), .Z1_t (new_AGEMA_signal_2052), .Z1_f (new_AGEMA_signal_2053) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (stateFF_MUX_inputPar_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_2051), .B1_t (new_AGEMA_signal_2052), .B1_f (new_AGEMA_signal_2053), .Z0_t (stateFF_MUX_inputPar_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_2910), .Z1_t (new_AGEMA_signal_2911), .Z1_f (new_AGEMA_signal_2912) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) stateFF_MUX_inputPar_mux_inst_63_U1_XOR2_U1 ( .A0_t (stateFF_MUX_inputPar_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_2910), .A1_t (new_AGEMA_signal_2911), .A1_f (new_AGEMA_signal_2912), .B0_t (data_out_s0_t[63]), .B0_f (data_out_s0_f[63]), .B1_t (data_out_s1_t[63]), .B1_f (data_out_s1_f[63]), .Z0_t (stateFF_inputPar[63]), .Z0_f (new_AGEMA_signal_3370), .Z1_t (new_AGEMA_signal_3371), .Z1_f (new_AGEMA_signal_3372) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U5 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (counter[3]), .A1_f (new_AGEMA_signal_1470), .B0_t (keyFF_outputPar[21]), .B0_f (new_AGEMA_signal_2054), .B1_t (new_AGEMA_signal_2055), .B1_f (new_AGEMA_signal_2056), .Z0_t (keyFF_counterAdd[3]), .Z0_f (new_AGEMA_signal_2057), .Z1_t (new_AGEMA_signal_2058), .Z1_f (new_AGEMA_signal_2059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U4 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (counter[1]), .A1_f (new_AGEMA_signal_1476), .B0_t (keyFF_outputPar[19]), .B0_f (new_AGEMA_signal_2060), .B1_t (new_AGEMA_signal_2061), .B1_f (new_AGEMA_signal_2062), .Z0_t (keyFF_counterAdd[1]), .Z0_f (new_AGEMA_signal_2063), .Z1_t (new_AGEMA_signal_2064), .Z1_f (new_AGEMA_signal_2065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U3 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (counter[4]), .A1_f (new_AGEMA_signal_1473), .B0_t (keyFF_outputPar[22]), .B0_f (new_AGEMA_signal_2066), .B1_t (new_AGEMA_signal_2067), .B1_f (new_AGEMA_signal_2068), .Z0_t (keyFF_counterAdd[4]), .Z0_f (new_AGEMA_signal_2069), .Z1_t (new_AGEMA_signal_2070), .Z1_f (new_AGEMA_signal_2071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U2 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (counter[0]), .A1_f (new_AGEMA_signal_1474), .B0_t (keyFF_outputPar[18]), .B0_f (new_AGEMA_signal_2072), .B1_t (new_AGEMA_signal_2073), .B1_f (new_AGEMA_signal_2074), .Z0_t (keyFF_counterAdd[0]), .Z0_f (new_AGEMA_signal_2075), .Z1_t (new_AGEMA_signal_2076), .Z1_f (new_AGEMA_signal_2077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (counter[2]), .A1_f (new_AGEMA_signal_1477), .B0_t (keyFF_outputPar[20]), .B0_f (new_AGEMA_signal_2078), .B1_t (new_AGEMA_signal_2079), .B1_f (new_AGEMA_signal_2080), .Z0_t (keyFF_counterAdd[2]), .Z0_f (new_AGEMA_signal_2081), .Z1_t (new_AGEMA_signal_2082), .Z1_f (new_AGEMA_signal_2083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (roundkey[0]), .A0_f (new_AGEMA_signal_1452), .A1_t (new_AGEMA_signal_1453), .A1_f (new_AGEMA_signal_1454), .B0_t (keyFF_inputPar[0]), .B0_f (new_AGEMA_signal_3373), .B1_t (new_AGEMA_signal_3374), .B1_f (new_AGEMA_signal_3375), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3797), .Z1_t (new_AGEMA_signal_3798), .Z1_f (new_AGEMA_signal_3799) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3797), .B1_t (new_AGEMA_signal_3798), .B1_f (new_AGEMA_signal_3799), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4219), .Z1_t (new_AGEMA_signal_4220), .Z1_f (new_AGEMA_signal_4221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4219), .A1_t (new_AGEMA_signal_4220), .A1_f (new_AGEMA_signal_4221), .B0_t (roundkey[0]), .B0_f (new_AGEMA_signal_1452), .B1_t (new_AGEMA_signal_1453), .B1_f (new_AGEMA_signal_1454), .Z0_t (keyRegKS[1]), .Z0_f (new_AGEMA_signal_3159), .Z1_t (new_AGEMA_signal_3160), .Z1_f (new_AGEMA_signal_3161) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (roundkey[1]), .A0_f (new_AGEMA_signal_1434), .A1_t (new_AGEMA_signal_1435), .A1_f (new_AGEMA_signal_1436), .B0_t (keyFF_inputPar[1]), .B0_f (new_AGEMA_signal_3376), .B1_t (new_AGEMA_signal_3377), .B1_f (new_AGEMA_signal_3378), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3800), .Z1_t (new_AGEMA_signal_3801), .Z1_f (new_AGEMA_signal_3802) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3800), .B1_t (new_AGEMA_signal_3801), .B1_f (new_AGEMA_signal_3802), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4222), .Z1_t (new_AGEMA_signal_4223), .Z1_f (new_AGEMA_signal_4224) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4222), .A1_t (new_AGEMA_signal_4223), .A1_f (new_AGEMA_signal_4224), .B0_t (roundkey[1]), .B0_f (new_AGEMA_signal_1434), .B1_t (new_AGEMA_signal_1435), .B1_f (new_AGEMA_signal_1436), .Z0_t (keyRegKS[2]), .Z0_f (new_AGEMA_signal_3165), .Z1_t (new_AGEMA_signal_3166), .Z1_f (new_AGEMA_signal_3167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (roundkey[2]), .A0_f (new_AGEMA_signal_1443), .A1_t (new_AGEMA_signal_1444), .A1_f (new_AGEMA_signal_1445), .B0_t (keyFF_inputPar[2]), .B0_f (new_AGEMA_signal_3379), .B1_t (new_AGEMA_signal_3380), .B1_f (new_AGEMA_signal_3381), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3803), .Z1_t (new_AGEMA_signal_3804), .Z1_f (new_AGEMA_signal_3805) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3803), .B1_t (new_AGEMA_signal_3804), .B1_f (new_AGEMA_signal_3805), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4225), .Z1_t (new_AGEMA_signal_4226), .Z1_f (new_AGEMA_signal_4227) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4225), .A1_t (new_AGEMA_signal_4226), .A1_f (new_AGEMA_signal_4227), .B0_t (roundkey[2]), .B0_f (new_AGEMA_signal_1443), .B1_t (new_AGEMA_signal_1444), .B1_f (new_AGEMA_signal_1445), .Z0_t (keyRegKS[3]), .Z0_f (new_AGEMA_signal_3171), .Z1_t (new_AGEMA_signal_3172), .Z1_f (new_AGEMA_signal_3173) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (roundkey[3]), .A0_f (new_AGEMA_signal_1461), .A1_t (new_AGEMA_signal_1462), .A1_f (new_AGEMA_signal_1463), .B0_t (keyFF_inputPar[3]), .B0_f (new_AGEMA_signal_3382), .B1_t (new_AGEMA_signal_3383), .B1_f (new_AGEMA_signal_3384), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3806), .Z1_t (new_AGEMA_signal_3807), .Z1_f (new_AGEMA_signal_3808) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3806), .B1_t (new_AGEMA_signal_3807), .B1_f (new_AGEMA_signal_3808), .Z0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4228), .Z1_t (new_AGEMA_signal_4229), .Z1_f (new_AGEMA_signal_4230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4228), .A1_t (new_AGEMA_signal_4229), .A1_f (new_AGEMA_signal_4230), .B0_t (roundkey[3]), .B0_f (new_AGEMA_signal_1461), .B1_t (new_AGEMA_signal_1462), .B1_f (new_AGEMA_signal_1463), .Z0_t (keyFF_outputPar[3]), .Z0_f (new_AGEMA_signal_2084), .Z1_t (new_AGEMA_signal_2085), .Z1_f (new_AGEMA_signal_2086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyRegKS[1]), .A0_f (new_AGEMA_signal_3159), .A1_t (new_AGEMA_signal_3160), .A1_f (new_AGEMA_signal_3161), .B0_t (keyFF_inputPar[4]), .B0_f (new_AGEMA_signal_3385), .B1_t (new_AGEMA_signal_3386), .B1_f (new_AGEMA_signal_3387), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3809), .Z1_t (new_AGEMA_signal_3810), .Z1_f (new_AGEMA_signal_3811) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3809), .B1_t (new_AGEMA_signal_3810), .B1_f (new_AGEMA_signal_3811), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4231), .Z1_t (new_AGEMA_signal_4232), .Z1_f (new_AGEMA_signal_4233) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4231), .A1_t (new_AGEMA_signal_4232), .A1_f (new_AGEMA_signal_4233), .B0_t (keyRegKS[1]), .B0_f (new_AGEMA_signal_3159), .B1_t (new_AGEMA_signal_3160), .B1_f (new_AGEMA_signal_3161), .Z0_t (keyFF_outputPar[4]), .Z0_f (new_AGEMA_signal_2093), .Z1_t (new_AGEMA_signal_2094), .Z1_f (new_AGEMA_signal_2095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyRegKS[2]), .A0_f (new_AGEMA_signal_3165), .A1_t (new_AGEMA_signal_3166), .A1_f (new_AGEMA_signal_3167), .B0_t (keyFF_inputPar[5]), .B0_f (new_AGEMA_signal_3388), .B1_t (new_AGEMA_signal_3389), .B1_f (new_AGEMA_signal_3390), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3812), .Z1_t (new_AGEMA_signal_3813), .Z1_f (new_AGEMA_signal_3814) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3812), .B1_t (new_AGEMA_signal_3813), .B1_f (new_AGEMA_signal_3814), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4234), .Z1_t (new_AGEMA_signal_4235), .Z1_f (new_AGEMA_signal_4236) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4234), .A1_t (new_AGEMA_signal_4235), .A1_f (new_AGEMA_signal_4236), .B0_t (keyRegKS[2]), .B0_f (new_AGEMA_signal_3165), .B1_t (new_AGEMA_signal_3166), .B1_f (new_AGEMA_signal_3167), .Z0_t (keyFF_outputPar[5]), .Z0_f (new_AGEMA_signal_2102), .Z1_t (new_AGEMA_signal_2103), .Z1_f (new_AGEMA_signal_2104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyRegKS[3]), .A0_f (new_AGEMA_signal_3171), .A1_t (new_AGEMA_signal_3172), .A1_f (new_AGEMA_signal_3173), .B0_t (keyFF_inputPar[6]), .B0_f (new_AGEMA_signal_3391), .B1_t (new_AGEMA_signal_3392), .B1_f (new_AGEMA_signal_3393), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3815), .Z1_t (new_AGEMA_signal_3816), .Z1_f (new_AGEMA_signal_3817) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3815), .B1_t (new_AGEMA_signal_3816), .B1_f (new_AGEMA_signal_3817), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4237), .Z1_t (new_AGEMA_signal_4238), .Z1_f (new_AGEMA_signal_4239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4237), .A1_t (new_AGEMA_signal_4238), .A1_f (new_AGEMA_signal_4239), .B0_t (keyRegKS[3]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (keyFF_outputPar[6]), .Z0_f (new_AGEMA_signal_2111), .Z1_t (new_AGEMA_signal_2112), .Z1_f (new_AGEMA_signal_2113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[3]), .A0_f (new_AGEMA_signal_2084), .A1_t (new_AGEMA_signal_2085), .A1_f (new_AGEMA_signal_2086), .B0_t (keyFF_inputPar[7]), .B0_f (new_AGEMA_signal_3394), .B1_t (new_AGEMA_signal_3395), .B1_f (new_AGEMA_signal_3396), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3818), .Z1_t (new_AGEMA_signal_3819), .Z1_f (new_AGEMA_signal_3820) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3818), .B1_t (new_AGEMA_signal_3819), .B1_f (new_AGEMA_signal_3820), .Z0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4240), .Z1_t (new_AGEMA_signal_4241), .Z1_f (new_AGEMA_signal_4242) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4240), .A1_t (new_AGEMA_signal_4241), .A1_f (new_AGEMA_signal_4242), .B0_t (keyFF_outputPar[3]), .B0_f (new_AGEMA_signal_2084), .B1_t (new_AGEMA_signal_2085), .B1_f (new_AGEMA_signal_2086), .Z0_t (keyFF_outputPar[7]), .Z0_f (new_AGEMA_signal_2120), .Z1_t (new_AGEMA_signal_2121), .Z1_f (new_AGEMA_signal_2122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[4]), .A0_f (new_AGEMA_signal_2093), .A1_t (new_AGEMA_signal_2094), .A1_f (new_AGEMA_signal_2095), .B0_t (keyFF_inputPar[8]), .B0_f (new_AGEMA_signal_3397), .B1_t (new_AGEMA_signal_3398), .B1_f (new_AGEMA_signal_3399), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3821), .Z1_t (new_AGEMA_signal_3822), .Z1_f (new_AGEMA_signal_3823) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3821), .B1_t (new_AGEMA_signal_3822), .B1_f (new_AGEMA_signal_3823), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4243), .Z1_t (new_AGEMA_signal_4244), .Z1_f (new_AGEMA_signal_4245) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4243), .A1_t (new_AGEMA_signal_4244), .A1_f (new_AGEMA_signal_4245), .B0_t (keyFF_outputPar[4]), .B0_f (new_AGEMA_signal_2093), .B1_t (new_AGEMA_signal_2094), .B1_f (new_AGEMA_signal_2095), .Z0_t (keyFF_outputPar[8]), .Z0_f (new_AGEMA_signal_2129), .Z1_t (new_AGEMA_signal_2130), .Z1_f (new_AGEMA_signal_2131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[5]), .A0_f (new_AGEMA_signal_2102), .A1_t (new_AGEMA_signal_2103), .A1_f (new_AGEMA_signal_2104), .B0_t (keyFF_inputPar[9]), .B0_f (new_AGEMA_signal_3400), .B1_t (new_AGEMA_signal_3401), .B1_f (new_AGEMA_signal_3402), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3824), .Z1_t (new_AGEMA_signal_3825), .Z1_f (new_AGEMA_signal_3826) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3824), .B1_t (new_AGEMA_signal_3825), .B1_f (new_AGEMA_signal_3826), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4246), .Z1_t (new_AGEMA_signal_4247), .Z1_f (new_AGEMA_signal_4248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4246), .A1_t (new_AGEMA_signal_4247), .A1_f (new_AGEMA_signal_4248), .B0_t (keyFF_outputPar[5]), .B0_f (new_AGEMA_signal_2102), .B1_t (new_AGEMA_signal_2103), .B1_f (new_AGEMA_signal_2104), .Z0_t (keyFF_outputPar[9]), .Z0_f (new_AGEMA_signal_2138), .Z1_t (new_AGEMA_signal_2139), .Z1_f (new_AGEMA_signal_2140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[6]), .A0_f (new_AGEMA_signal_2111), .A1_t (new_AGEMA_signal_2112), .A1_f (new_AGEMA_signal_2113), .B0_t (keyFF_inputPar[10]), .B0_f (new_AGEMA_signal_3403), .B1_t (new_AGEMA_signal_3404), .B1_f (new_AGEMA_signal_3405), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3827), .Z1_t (new_AGEMA_signal_3828), .Z1_f (new_AGEMA_signal_3829) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3827), .B1_t (new_AGEMA_signal_3828), .B1_f (new_AGEMA_signal_3829), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4249), .Z1_t (new_AGEMA_signal_4250), .Z1_f (new_AGEMA_signal_4251) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4249), .A1_t (new_AGEMA_signal_4250), .A1_f (new_AGEMA_signal_4251), .B0_t (keyFF_outputPar[6]), .B0_f (new_AGEMA_signal_2111), .B1_t (new_AGEMA_signal_2112), .B1_f (new_AGEMA_signal_2113), .Z0_t (keyFF_outputPar[10]), .Z0_f (new_AGEMA_signal_2147), .Z1_t (new_AGEMA_signal_2148), .Z1_f (new_AGEMA_signal_2149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[7]), .A0_f (new_AGEMA_signal_2120), .A1_t (new_AGEMA_signal_2121), .A1_f (new_AGEMA_signal_2122), .B0_t (keyFF_inputPar[11]), .B0_f (new_AGEMA_signal_3406), .B1_t (new_AGEMA_signal_3407), .B1_f (new_AGEMA_signal_3408), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3830), .Z1_t (new_AGEMA_signal_3831), .Z1_f (new_AGEMA_signal_3832) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3830), .B1_t (new_AGEMA_signal_3831), .B1_f (new_AGEMA_signal_3832), .Z0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4252), .Z1_t (new_AGEMA_signal_4253), .Z1_f (new_AGEMA_signal_4254) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4252), .A1_t (new_AGEMA_signal_4253), .A1_f (new_AGEMA_signal_4254), .B0_t (keyFF_outputPar[7]), .B0_f (new_AGEMA_signal_2120), .B1_t (new_AGEMA_signal_2121), .B1_f (new_AGEMA_signal_2122), .Z0_t (keyFF_outputPar[11]), .Z0_f (new_AGEMA_signal_2156), .Z1_t (new_AGEMA_signal_2157), .Z1_f (new_AGEMA_signal_2158) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[8]), .A0_f (new_AGEMA_signal_2129), .A1_t (new_AGEMA_signal_2130), .A1_f (new_AGEMA_signal_2131), .B0_t (keyFF_inputPar[12]), .B0_f (new_AGEMA_signal_3409), .B1_t (new_AGEMA_signal_3410), .B1_f (new_AGEMA_signal_3411), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3833), .Z1_t (new_AGEMA_signal_3834), .Z1_f (new_AGEMA_signal_3835) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3833), .B1_t (new_AGEMA_signal_3834), .B1_f (new_AGEMA_signal_3835), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4255), .Z1_t (new_AGEMA_signal_4256), .Z1_f (new_AGEMA_signal_4257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4255), .A1_t (new_AGEMA_signal_4256), .A1_f (new_AGEMA_signal_4257), .B0_t (keyFF_outputPar[8]), .B0_f (new_AGEMA_signal_2129), .B1_t (new_AGEMA_signal_2130), .B1_f (new_AGEMA_signal_2131), .Z0_t (keyFF_outputPar[12]), .Z0_f (new_AGEMA_signal_2165), .Z1_t (new_AGEMA_signal_2166), .Z1_f (new_AGEMA_signal_2167) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[9]), .A0_f (new_AGEMA_signal_2138), .A1_t (new_AGEMA_signal_2139), .A1_f (new_AGEMA_signal_2140), .B0_t (keyFF_inputPar[13]), .B0_f (new_AGEMA_signal_3412), .B1_t (new_AGEMA_signal_3413), .B1_f (new_AGEMA_signal_3414), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3836), .Z1_t (new_AGEMA_signal_3837), .Z1_f (new_AGEMA_signal_3838) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3836), .B1_t (new_AGEMA_signal_3837), .B1_f (new_AGEMA_signal_3838), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4258), .Z1_t (new_AGEMA_signal_4259), .Z1_f (new_AGEMA_signal_4260) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4258), .A1_t (new_AGEMA_signal_4259), .A1_f (new_AGEMA_signal_4260), .B0_t (keyFF_outputPar[9]), .B0_f (new_AGEMA_signal_2138), .B1_t (new_AGEMA_signal_2139), .B1_f (new_AGEMA_signal_2140), .Z0_t (keyFF_outputPar[13]), .Z0_f (new_AGEMA_signal_2174), .Z1_t (new_AGEMA_signal_2175), .Z1_f (new_AGEMA_signal_2176) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[10]), .A0_f (new_AGEMA_signal_2147), .A1_t (new_AGEMA_signal_2148), .A1_f (new_AGEMA_signal_2149), .B0_t (keyFF_inputPar[14]), .B0_f (new_AGEMA_signal_3415), .B1_t (new_AGEMA_signal_3416), .B1_f (new_AGEMA_signal_3417), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3839), .Z1_t (new_AGEMA_signal_3840), .Z1_f (new_AGEMA_signal_3841) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3839), .B1_t (new_AGEMA_signal_3840), .B1_f (new_AGEMA_signal_3841), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4261), .Z1_t (new_AGEMA_signal_4262), .Z1_f (new_AGEMA_signal_4263) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4261), .A1_t (new_AGEMA_signal_4262), .A1_f (new_AGEMA_signal_4263), .B0_t (keyFF_outputPar[10]), .B0_f (new_AGEMA_signal_2147), .B1_t (new_AGEMA_signal_2148), .B1_f (new_AGEMA_signal_2149), .Z0_t (keyFF_outputPar[14]), .Z0_f (new_AGEMA_signal_2183), .Z1_t (new_AGEMA_signal_2184), .Z1_f (new_AGEMA_signal_2185) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[11]), .A0_f (new_AGEMA_signal_2156), .A1_t (new_AGEMA_signal_2157), .A1_f (new_AGEMA_signal_2158), .B0_t (keyFF_inputPar[15]), .B0_f (new_AGEMA_signal_4010), .B1_t (new_AGEMA_signal_4011), .B1_f (new_AGEMA_signal_4012), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4264), .Z1_t (new_AGEMA_signal_4265), .Z1_f (new_AGEMA_signal_4266) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4264), .B1_t (new_AGEMA_signal_4265), .B1_f (new_AGEMA_signal_4266), .Z0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4464), .Z1_t (new_AGEMA_signal_4465), .Z1_f (new_AGEMA_signal_4466) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4464), .A1_t (new_AGEMA_signal_4465), .A1_f (new_AGEMA_signal_4466), .B0_t (keyFF_outputPar[11]), .B0_f (new_AGEMA_signal_2156), .B1_t (new_AGEMA_signal_2157), .B1_f (new_AGEMA_signal_2158), .Z0_t (keyFF_outputPar[15]), .Z0_f (new_AGEMA_signal_2192), .Z1_t (new_AGEMA_signal_2193), .Z1_f (new_AGEMA_signal_2194) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[12]), .A0_f (new_AGEMA_signal_2165), .A1_t (new_AGEMA_signal_2166), .A1_f (new_AGEMA_signal_2167), .B0_t (keyFF_inputPar[16]), .B0_f (new_AGEMA_signal_4013), .B1_t (new_AGEMA_signal_4014), .B1_f (new_AGEMA_signal_4015), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_4267), .Z1_t (new_AGEMA_signal_4268), .Z1_f (new_AGEMA_signal_4269) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_4267), .B1_t (new_AGEMA_signal_4268), .B1_f (new_AGEMA_signal_4269), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4467), .Z1_t (new_AGEMA_signal_4468), .Z1_f (new_AGEMA_signal_4469) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4467), .A1_t (new_AGEMA_signal_4468), .A1_f (new_AGEMA_signal_4469), .B0_t (keyFF_outputPar[12]), .B0_f (new_AGEMA_signal_2165), .B1_t (new_AGEMA_signal_2166), .B1_f (new_AGEMA_signal_2167), .Z0_t (keyFF_outputPar[16]), .Z0_f (new_AGEMA_signal_2201), .Z1_t (new_AGEMA_signal_2202), .Z1_f (new_AGEMA_signal_2203) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[13]), .A0_f (new_AGEMA_signal_2174), .A1_t (new_AGEMA_signal_2175), .A1_f (new_AGEMA_signal_2176), .B0_t (keyFF_inputPar[17]), .B0_f (new_AGEMA_signal_4016), .B1_t (new_AGEMA_signal_4017), .B1_f (new_AGEMA_signal_4018), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4270), .Z1_t (new_AGEMA_signal_4271), .Z1_f (new_AGEMA_signal_4272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4270), .B1_t (new_AGEMA_signal_4271), .B1_f (new_AGEMA_signal_4272), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4470), .Z1_t (new_AGEMA_signal_4471), .Z1_f (new_AGEMA_signal_4472) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4470), .A1_t (new_AGEMA_signal_4471), .A1_f (new_AGEMA_signal_4472), .B0_t (keyFF_outputPar[13]), .B0_f (new_AGEMA_signal_2174), .B1_t (new_AGEMA_signal_2175), .B1_f (new_AGEMA_signal_2176), .Z0_t (keyFF_outputPar[17]), .Z0_f (new_AGEMA_signal_2210), .Z1_t (new_AGEMA_signal_2211), .Z1_f (new_AGEMA_signal_2212) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[14]), .A0_f (new_AGEMA_signal_2183), .A1_t (new_AGEMA_signal_2184), .A1_f (new_AGEMA_signal_2185), .B0_t (keyFF_inputPar[18]), .B0_f (new_AGEMA_signal_4019), .B1_t (new_AGEMA_signal_4020), .B1_f (new_AGEMA_signal_4021), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_4273), .Z1_t (new_AGEMA_signal_4274), .Z1_f (new_AGEMA_signal_4275) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_4273), .B1_t (new_AGEMA_signal_4274), .B1_f (new_AGEMA_signal_4275), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4473), .Z1_t (new_AGEMA_signal_4474), .Z1_f (new_AGEMA_signal_4475) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4473), .A1_t (new_AGEMA_signal_4474), .A1_f (new_AGEMA_signal_4475), .B0_t (keyFF_outputPar[14]), .B0_f (new_AGEMA_signal_2183), .B1_t (new_AGEMA_signal_2184), .B1_f (new_AGEMA_signal_2185), .Z0_t (keyFF_outputPar[18]), .Z0_f (new_AGEMA_signal_2072), .Z1_t (new_AGEMA_signal_2073), .Z1_f (new_AGEMA_signal_2074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[15]), .A0_f (new_AGEMA_signal_2192), .A1_t (new_AGEMA_signal_2193), .A1_f (new_AGEMA_signal_2194), .B0_t (keyFF_inputPar[19]), .B0_f (new_AGEMA_signal_4022), .B1_t (new_AGEMA_signal_4023), .B1_f (new_AGEMA_signal_4024), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4276), .Z1_t (new_AGEMA_signal_4277), .Z1_f (new_AGEMA_signal_4278) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4276), .B1_t (new_AGEMA_signal_4277), .B1_f (new_AGEMA_signal_4278), .Z0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4476), .Z1_t (new_AGEMA_signal_4477), .Z1_f (new_AGEMA_signal_4478) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4476), .A1_t (new_AGEMA_signal_4477), .A1_f (new_AGEMA_signal_4478), .B0_t (keyFF_outputPar[15]), .B0_f (new_AGEMA_signal_2192), .B1_t (new_AGEMA_signal_2193), .B1_f (new_AGEMA_signal_2194), .Z0_t (keyFF_outputPar[19]), .Z0_f (new_AGEMA_signal_2060), .Z1_t (new_AGEMA_signal_2061), .Z1_f (new_AGEMA_signal_2062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[16]), .A0_f (new_AGEMA_signal_2201), .A1_t (new_AGEMA_signal_2202), .A1_f (new_AGEMA_signal_2203), .B0_t (keyFF_inputPar[20]), .B0_f (new_AGEMA_signal_3433), .B1_t (new_AGEMA_signal_3434), .B1_f (new_AGEMA_signal_3435), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3842), .Z1_t (new_AGEMA_signal_3843), .Z1_f (new_AGEMA_signal_3844) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3842), .B1_t (new_AGEMA_signal_3843), .B1_f (new_AGEMA_signal_3844), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4279), .Z1_t (new_AGEMA_signal_4280), .Z1_f (new_AGEMA_signal_4281) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4279), .A1_t (new_AGEMA_signal_4280), .A1_f (new_AGEMA_signal_4281), .B0_t (keyFF_outputPar[16]), .B0_f (new_AGEMA_signal_2201), .B1_t (new_AGEMA_signal_2202), .B1_f (new_AGEMA_signal_2203), .Z0_t (keyFF_outputPar[20]), .Z0_f (new_AGEMA_signal_2078), .Z1_t (new_AGEMA_signal_2079), .Z1_f (new_AGEMA_signal_2080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[17]), .A0_f (new_AGEMA_signal_2210), .A1_t (new_AGEMA_signal_2211), .A1_f (new_AGEMA_signal_2212), .B0_t (keyFF_inputPar[21]), .B0_f (new_AGEMA_signal_3436), .B1_t (new_AGEMA_signal_3437), .B1_f (new_AGEMA_signal_3438), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3845), .Z1_t (new_AGEMA_signal_3846), .Z1_f (new_AGEMA_signal_3847) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3845), .B1_t (new_AGEMA_signal_3846), .B1_f (new_AGEMA_signal_3847), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4282), .Z1_t (new_AGEMA_signal_4283), .Z1_f (new_AGEMA_signal_4284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4282), .A1_t (new_AGEMA_signal_4283), .A1_f (new_AGEMA_signal_4284), .B0_t (keyFF_outputPar[17]), .B0_f (new_AGEMA_signal_2210), .B1_t (new_AGEMA_signal_2211), .B1_f (new_AGEMA_signal_2212), .Z0_t (keyFF_outputPar[21]), .Z0_f (new_AGEMA_signal_2054), .Z1_t (new_AGEMA_signal_2055), .Z1_f (new_AGEMA_signal_2056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[18]), .A0_f (new_AGEMA_signal_2072), .A1_t (new_AGEMA_signal_2073), .A1_f (new_AGEMA_signal_2074), .B0_t (keyFF_inputPar[22]), .B0_f (new_AGEMA_signal_3439), .B1_t (new_AGEMA_signal_3440), .B1_f (new_AGEMA_signal_3441), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3848), .Z1_t (new_AGEMA_signal_3849), .Z1_f (new_AGEMA_signal_3850) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3848), .B1_t (new_AGEMA_signal_3849), .B1_f (new_AGEMA_signal_3850), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4285), .Z1_t (new_AGEMA_signal_4286), .Z1_f (new_AGEMA_signal_4287) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4285), .A1_t (new_AGEMA_signal_4286), .A1_f (new_AGEMA_signal_4287), .B0_t (keyFF_outputPar[18]), .B0_f (new_AGEMA_signal_2072), .B1_t (new_AGEMA_signal_2073), .B1_f (new_AGEMA_signal_2074), .Z0_t (keyFF_outputPar[22]), .Z0_f (new_AGEMA_signal_2066), .Z1_t (new_AGEMA_signal_2067), .Z1_f (new_AGEMA_signal_2068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[19]), .A0_f (new_AGEMA_signal_2060), .A1_t (new_AGEMA_signal_2061), .A1_f (new_AGEMA_signal_2062), .B0_t (keyFF_inputPar[23]), .B0_f (new_AGEMA_signal_3442), .B1_t (new_AGEMA_signal_3443), .B1_f (new_AGEMA_signal_3444), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3851), .Z1_t (new_AGEMA_signal_3852), .Z1_f (new_AGEMA_signal_3853) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3851), .B1_t (new_AGEMA_signal_3852), .B1_f (new_AGEMA_signal_3853), .Z0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4288), .Z1_t (new_AGEMA_signal_4289), .Z1_f (new_AGEMA_signal_4290) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4288), .A1_t (new_AGEMA_signal_4289), .A1_f (new_AGEMA_signal_4290), .B0_t (keyFF_outputPar[19]), .B0_f (new_AGEMA_signal_2060), .B1_t (new_AGEMA_signal_2061), .B1_f (new_AGEMA_signal_2062), .Z0_t (keyFF_outputPar[23]), .Z0_f (new_AGEMA_signal_2219), .Z1_t (new_AGEMA_signal_2220), .Z1_f (new_AGEMA_signal_2221) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[20]), .A0_f (new_AGEMA_signal_2078), .A1_t (new_AGEMA_signal_2079), .A1_f (new_AGEMA_signal_2080), .B0_t (keyFF_inputPar[24]), .B0_f (new_AGEMA_signal_3445), .B1_t (new_AGEMA_signal_3446), .B1_f (new_AGEMA_signal_3447), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3854), .Z1_t (new_AGEMA_signal_3855), .Z1_f (new_AGEMA_signal_3856) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3854), .B1_t (new_AGEMA_signal_3855), .B1_f (new_AGEMA_signal_3856), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4291), .Z1_t (new_AGEMA_signal_4292), .Z1_f (new_AGEMA_signal_4293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4291), .A1_t (new_AGEMA_signal_4292), .A1_f (new_AGEMA_signal_4293), .B0_t (keyFF_outputPar[20]), .B0_f (new_AGEMA_signal_2078), .B1_t (new_AGEMA_signal_2079), .B1_f (new_AGEMA_signal_2080), .Z0_t (keyFF_outputPar[24]), .Z0_f (new_AGEMA_signal_2228), .Z1_t (new_AGEMA_signal_2229), .Z1_f (new_AGEMA_signal_2230) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[21]), .A0_f (new_AGEMA_signal_2054), .A1_t (new_AGEMA_signal_2055), .A1_f (new_AGEMA_signal_2056), .B0_t (keyFF_inputPar[25]), .B0_f (new_AGEMA_signal_3448), .B1_t (new_AGEMA_signal_3449), .B1_f (new_AGEMA_signal_3450), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3857), .Z1_t (new_AGEMA_signal_3858), .Z1_f (new_AGEMA_signal_3859) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3857), .B1_t (new_AGEMA_signal_3858), .B1_f (new_AGEMA_signal_3859), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4294), .Z1_t (new_AGEMA_signal_4295), .Z1_f (new_AGEMA_signal_4296) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4294), .A1_t (new_AGEMA_signal_4295), .A1_f (new_AGEMA_signal_4296), .B0_t (keyFF_outputPar[21]), .B0_f (new_AGEMA_signal_2054), .B1_t (new_AGEMA_signal_2055), .B1_f (new_AGEMA_signal_2056), .Z0_t (keyFF_outputPar[25]), .Z0_f (new_AGEMA_signal_2237), .Z1_t (new_AGEMA_signal_2238), .Z1_f (new_AGEMA_signal_2239) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[22]), .A0_f (new_AGEMA_signal_2066), .A1_t (new_AGEMA_signal_2067), .A1_f (new_AGEMA_signal_2068), .B0_t (keyFF_inputPar[26]), .B0_f (new_AGEMA_signal_3451), .B1_t (new_AGEMA_signal_3452), .B1_f (new_AGEMA_signal_3453), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3860), .Z1_t (new_AGEMA_signal_3861), .Z1_f (new_AGEMA_signal_3862) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3860), .B1_t (new_AGEMA_signal_3861), .B1_f (new_AGEMA_signal_3862), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4297), .Z1_t (new_AGEMA_signal_4298), .Z1_f (new_AGEMA_signal_4299) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4297), .A1_t (new_AGEMA_signal_4298), .A1_f (new_AGEMA_signal_4299), .B0_t (keyFF_outputPar[22]), .B0_f (new_AGEMA_signal_2066), .B1_t (new_AGEMA_signal_2067), .B1_f (new_AGEMA_signal_2068), .Z0_t (keyFF_outputPar[26]), .Z0_f (new_AGEMA_signal_2246), .Z1_t (new_AGEMA_signal_2247), .Z1_f (new_AGEMA_signal_2248) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[23]), .A0_f (new_AGEMA_signal_2219), .A1_t (new_AGEMA_signal_2220), .A1_f (new_AGEMA_signal_2221), .B0_t (keyFF_inputPar[27]), .B0_f (new_AGEMA_signal_3454), .B1_t (new_AGEMA_signal_3455), .B1_f (new_AGEMA_signal_3456), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3863), .Z1_t (new_AGEMA_signal_3864), .Z1_f (new_AGEMA_signal_3865) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3863), .B1_t (new_AGEMA_signal_3864), .B1_f (new_AGEMA_signal_3865), .Z0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4300), .Z1_t (new_AGEMA_signal_4301), .Z1_f (new_AGEMA_signal_4302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4300), .A1_t (new_AGEMA_signal_4301), .A1_f (new_AGEMA_signal_4302), .B0_t (keyFF_outputPar[23]), .B0_f (new_AGEMA_signal_2219), .B1_t (new_AGEMA_signal_2220), .B1_f (new_AGEMA_signal_2221), .Z0_t (keyFF_outputPar[27]), .Z0_f (new_AGEMA_signal_2255), .Z1_t (new_AGEMA_signal_2256), .Z1_f (new_AGEMA_signal_2257) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[24]), .A0_f (new_AGEMA_signal_2228), .A1_t (new_AGEMA_signal_2229), .A1_f (new_AGEMA_signal_2230), .B0_t (keyFF_inputPar[28]), .B0_f (new_AGEMA_signal_3457), .B1_t (new_AGEMA_signal_3458), .B1_f (new_AGEMA_signal_3459), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3866), .Z1_t (new_AGEMA_signal_3867), .Z1_f (new_AGEMA_signal_3868) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3866), .B1_t (new_AGEMA_signal_3867), .B1_f (new_AGEMA_signal_3868), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4303), .Z1_t (new_AGEMA_signal_4304), .Z1_f (new_AGEMA_signal_4305) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4303), .A1_t (new_AGEMA_signal_4304), .A1_f (new_AGEMA_signal_4305), .B0_t (keyFF_outputPar[24]), .B0_f (new_AGEMA_signal_2228), .B1_t (new_AGEMA_signal_2229), .B1_f (new_AGEMA_signal_2230), .Z0_t (keyFF_outputPar[28]), .Z0_f (new_AGEMA_signal_2264), .Z1_t (new_AGEMA_signal_2265), .Z1_f (new_AGEMA_signal_2266) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[25]), .A0_f (new_AGEMA_signal_2237), .A1_t (new_AGEMA_signal_2238), .A1_f (new_AGEMA_signal_2239), .B0_t (keyFF_inputPar[29]), .B0_f (new_AGEMA_signal_3460), .B1_t (new_AGEMA_signal_3461), .B1_f (new_AGEMA_signal_3462), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3869), .Z1_t (new_AGEMA_signal_3870), .Z1_f (new_AGEMA_signal_3871) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3869), .B1_t (new_AGEMA_signal_3870), .B1_f (new_AGEMA_signal_3871), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4306), .Z1_t (new_AGEMA_signal_4307), .Z1_f (new_AGEMA_signal_4308) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4306), .A1_t (new_AGEMA_signal_4307), .A1_f (new_AGEMA_signal_4308), .B0_t (keyFF_outputPar[25]), .B0_f (new_AGEMA_signal_2237), .B1_t (new_AGEMA_signal_2238), .B1_f (new_AGEMA_signal_2239), .Z0_t (keyFF_outputPar[29]), .Z0_f (new_AGEMA_signal_2273), .Z1_t (new_AGEMA_signal_2274), .Z1_f (new_AGEMA_signal_2275) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[26]), .A0_f (new_AGEMA_signal_2246), .A1_t (new_AGEMA_signal_2247), .A1_f (new_AGEMA_signal_2248), .B0_t (keyFF_inputPar[30]), .B0_f (new_AGEMA_signal_3463), .B1_t (new_AGEMA_signal_3464), .B1_f (new_AGEMA_signal_3465), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3872), .Z1_t (new_AGEMA_signal_3873), .Z1_f (new_AGEMA_signal_3874) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3872), .B1_t (new_AGEMA_signal_3873), .B1_f (new_AGEMA_signal_3874), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4309), .Z1_t (new_AGEMA_signal_4310), .Z1_f (new_AGEMA_signal_4311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4309), .A1_t (new_AGEMA_signal_4310), .A1_f (new_AGEMA_signal_4311), .B0_t (keyFF_outputPar[26]), .B0_f (new_AGEMA_signal_2246), .B1_t (new_AGEMA_signal_2247), .B1_f (new_AGEMA_signal_2248), .Z0_t (keyFF_outputPar[30]), .Z0_f (new_AGEMA_signal_2282), .Z1_t (new_AGEMA_signal_2283), .Z1_f (new_AGEMA_signal_2284) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[27]), .A0_f (new_AGEMA_signal_2255), .A1_t (new_AGEMA_signal_2256), .A1_f (new_AGEMA_signal_2257), .B0_t (keyFF_inputPar[31]), .B0_f (new_AGEMA_signal_3466), .B1_t (new_AGEMA_signal_3467), .B1_f (new_AGEMA_signal_3468), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3875), .Z1_t (new_AGEMA_signal_3876), .Z1_f (new_AGEMA_signal_3877) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3875), .B1_t (new_AGEMA_signal_3876), .B1_f (new_AGEMA_signal_3877), .Z0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4312), .Z1_t (new_AGEMA_signal_4313), .Z1_f (new_AGEMA_signal_4314) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4312), .A1_t (new_AGEMA_signal_4313), .A1_f (new_AGEMA_signal_4314), .B0_t (keyFF_outputPar[27]), .B0_f (new_AGEMA_signal_2255), .B1_t (new_AGEMA_signal_2256), .B1_f (new_AGEMA_signal_2257), .Z0_t (keyFF_outputPar[31]), .Z0_f (new_AGEMA_signal_2291), .Z1_t (new_AGEMA_signal_2292), .Z1_f (new_AGEMA_signal_2293) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[28]), .A0_f (new_AGEMA_signal_2264), .A1_t (new_AGEMA_signal_2265), .A1_f (new_AGEMA_signal_2266), .B0_t (keyFF_inputPar[32]), .B0_f (new_AGEMA_signal_3469), .B1_t (new_AGEMA_signal_3470), .B1_f (new_AGEMA_signal_3471), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3878), .Z1_t (new_AGEMA_signal_3879), .Z1_f (new_AGEMA_signal_3880) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3878), .B1_t (new_AGEMA_signal_3879), .B1_f (new_AGEMA_signal_3880), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4315), .Z1_t (new_AGEMA_signal_4316), .Z1_f (new_AGEMA_signal_4317) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4315), .A1_t (new_AGEMA_signal_4316), .A1_f (new_AGEMA_signal_4317), .B0_t (keyFF_outputPar[28]), .B0_f (new_AGEMA_signal_2264), .B1_t (new_AGEMA_signal_2265), .B1_f (new_AGEMA_signal_2266), .Z0_t (keyFF_outputPar[32]), .Z0_f (new_AGEMA_signal_2300), .Z1_t (new_AGEMA_signal_2301), .Z1_f (new_AGEMA_signal_2302) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[29]), .A0_f (new_AGEMA_signal_2273), .A1_t (new_AGEMA_signal_2274), .A1_f (new_AGEMA_signal_2275), .B0_t (keyFF_inputPar[33]), .B0_f (new_AGEMA_signal_3472), .B1_t (new_AGEMA_signal_3473), .B1_f (new_AGEMA_signal_3474), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3881), .Z1_t (new_AGEMA_signal_3882), .Z1_f (new_AGEMA_signal_3883) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3881), .B1_t (new_AGEMA_signal_3882), .B1_f (new_AGEMA_signal_3883), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4318), .Z1_t (new_AGEMA_signal_4319), .Z1_f (new_AGEMA_signal_4320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4318), .A1_t (new_AGEMA_signal_4319), .A1_f (new_AGEMA_signal_4320), .B0_t (keyFF_outputPar[29]), .B0_f (new_AGEMA_signal_2273), .B1_t (new_AGEMA_signal_2274), .B1_f (new_AGEMA_signal_2275), .Z0_t (keyFF_outputPar[33]), .Z0_f (new_AGEMA_signal_2309), .Z1_t (new_AGEMA_signal_2310), .Z1_f (new_AGEMA_signal_2311) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[30]), .A0_f (new_AGEMA_signal_2282), .A1_t (new_AGEMA_signal_2283), .A1_f (new_AGEMA_signal_2284), .B0_t (keyFF_inputPar[34]), .B0_f (new_AGEMA_signal_3475), .B1_t (new_AGEMA_signal_3476), .B1_f (new_AGEMA_signal_3477), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3884), .Z1_t (new_AGEMA_signal_3885), .Z1_f (new_AGEMA_signal_3886) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3884), .B1_t (new_AGEMA_signal_3885), .B1_f (new_AGEMA_signal_3886), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4321), .Z1_t (new_AGEMA_signal_4322), .Z1_f (new_AGEMA_signal_4323) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4321), .A1_t (new_AGEMA_signal_4322), .A1_f (new_AGEMA_signal_4323), .B0_t (keyFF_outputPar[30]), .B0_f (new_AGEMA_signal_2282), .B1_t (new_AGEMA_signal_2283), .B1_f (new_AGEMA_signal_2284), .Z0_t (keyFF_outputPar[34]), .Z0_f (new_AGEMA_signal_2318), .Z1_t (new_AGEMA_signal_2319), .Z1_f (new_AGEMA_signal_2320) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[31]), .A0_f (new_AGEMA_signal_2291), .A1_t (new_AGEMA_signal_2292), .A1_f (new_AGEMA_signal_2293), .B0_t (keyFF_inputPar[35]), .B0_f (new_AGEMA_signal_3478), .B1_t (new_AGEMA_signal_3479), .B1_f (new_AGEMA_signal_3480), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3887), .Z1_t (new_AGEMA_signal_3888), .Z1_f (new_AGEMA_signal_3889) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3887), .B1_t (new_AGEMA_signal_3888), .B1_f (new_AGEMA_signal_3889), .Z0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4324), .Z1_t (new_AGEMA_signal_4325), .Z1_f (new_AGEMA_signal_4326) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4324), .A1_t (new_AGEMA_signal_4325), .A1_f (new_AGEMA_signal_4326), .B0_t (keyFF_outputPar[31]), .B0_f (new_AGEMA_signal_2291), .B1_t (new_AGEMA_signal_2292), .B1_f (new_AGEMA_signal_2293), .Z0_t (keyFF_outputPar[35]), .Z0_f (new_AGEMA_signal_2327), .Z1_t (new_AGEMA_signal_2328), .Z1_f (new_AGEMA_signal_2329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[32]), .A0_f (new_AGEMA_signal_2300), .A1_t (new_AGEMA_signal_2301), .A1_f (new_AGEMA_signal_2302), .B0_t (keyFF_inputPar[36]), .B0_f (new_AGEMA_signal_3481), .B1_t (new_AGEMA_signal_3482), .B1_f (new_AGEMA_signal_3483), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3890), .Z1_t (new_AGEMA_signal_3891), .Z1_f (new_AGEMA_signal_3892) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3890), .B1_t (new_AGEMA_signal_3891), .B1_f (new_AGEMA_signal_3892), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4327), .Z1_t (new_AGEMA_signal_4328), .Z1_f (new_AGEMA_signal_4329) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4327), .A1_t (new_AGEMA_signal_4328), .A1_f (new_AGEMA_signal_4329), .B0_t (keyFF_outputPar[32]), .B0_f (new_AGEMA_signal_2300), .B1_t (new_AGEMA_signal_2301), .B1_f (new_AGEMA_signal_2302), .Z0_t (keyFF_outputPar[36]), .Z0_f (new_AGEMA_signal_2336), .Z1_t (new_AGEMA_signal_2337), .Z1_f (new_AGEMA_signal_2338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[33]), .A0_f (new_AGEMA_signal_2309), .A1_t (new_AGEMA_signal_2310), .A1_f (new_AGEMA_signal_2311), .B0_t (keyFF_inputPar[37]), .B0_f (new_AGEMA_signal_3484), .B1_t (new_AGEMA_signal_3485), .B1_f (new_AGEMA_signal_3486), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3893), .Z1_t (new_AGEMA_signal_3894), .Z1_f (new_AGEMA_signal_3895) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3893), .B1_t (new_AGEMA_signal_3894), .B1_f (new_AGEMA_signal_3895), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4330), .Z1_t (new_AGEMA_signal_4331), .Z1_f (new_AGEMA_signal_4332) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4330), .A1_t (new_AGEMA_signal_4331), .A1_f (new_AGEMA_signal_4332), .B0_t (keyFF_outputPar[33]), .B0_f (new_AGEMA_signal_2309), .B1_t (new_AGEMA_signal_2310), .B1_f (new_AGEMA_signal_2311), .Z0_t (keyFF_outputPar[37]), .Z0_f (new_AGEMA_signal_2345), .Z1_t (new_AGEMA_signal_2346), .Z1_f (new_AGEMA_signal_2347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[34]), .A0_f (new_AGEMA_signal_2318), .A1_t (new_AGEMA_signal_2319), .A1_f (new_AGEMA_signal_2320), .B0_t (keyFF_inputPar[38]), .B0_f (new_AGEMA_signal_3487), .B1_t (new_AGEMA_signal_3488), .B1_f (new_AGEMA_signal_3489), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3896), .Z1_t (new_AGEMA_signal_3897), .Z1_f (new_AGEMA_signal_3898) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3896), .B1_t (new_AGEMA_signal_3897), .B1_f (new_AGEMA_signal_3898), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4333), .Z1_t (new_AGEMA_signal_4334), .Z1_f (new_AGEMA_signal_4335) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4333), .A1_t (new_AGEMA_signal_4334), .A1_f (new_AGEMA_signal_4335), .B0_t (keyFF_outputPar[34]), .B0_f (new_AGEMA_signal_2318), .B1_t (new_AGEMA_signal_2319), .B1_f (new_AGEMA_signal_2320), .Z0_t (keyFF_outputPar[38]), .Z0_f (new_AGEMA_signal_2354), .Z1_t (new_AGEMA_signal_2355), .Z1_f (new_AGEMA_signal_2356) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[35]), .A0_f (new_AGEMA_signal_2327), .A1_t (new_AGEMA_signal_2328), .A1_f (new_AGEMA_signal_2329), .B0_t (keyFF_inputPar[39]), .B0_f (new_AGEMA_signal_3490), .B1_t (new_AGEMA_signal_3491), .B1_f (new_AGEMA_signal_3492), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3899), .Z1_t (new_AGEMA_signal_3900), .Z1_f (new_AGEMA_signal_3901) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3899), .B1_t (new_AGEMA_signal_3900), .B1_f (new_AGEMA_signal_3901), .Z0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4336), .Z1_t (new_AGEMA_signal_4337), .Z1_f (new_AGEMA_signal_4338) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4336), .A1_t (new_AGEMA_signal_4337), .A1_f (new_AGEMA_signal_4338), .B0_t (keyFF_outputPar[35]), .B0_f (new_AGEMA_signal_2327), .B1_t (new_AGEMA_signal_2328), .B1_f (new_AGEMA_signal_2329), .Z0_t (keyFF_outputPar[39]), .Z0_f (new_AGEMA_signal_2363), .Z1_t (new_AGEMA_signal_2364), .Z1_f (new_AGEMA_signal_2365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[36]), .A0_f (new_AGEMA_signal_2336), .A1_t (new_AGEMA_signal_2337), .A1_f (new_AGEMA_signal_2338), .B0_t (keyFF_inputPar[40]), .B0_f (new_AGEMA_signal_3493), .B1_t (new_AGEMA_signal_3494), .B1_f (new_AGEMA_signal_3495), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3902), .Z1_t (new_AGEMA_signal_3903), .Z1_f (new_AGEMA_signal_3904) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3902), .B1_t (new_AGEMA_signal_3903), .B1_f (new_AGEMA_signal_3904), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4339), .Z1_t (new_AGEMA_signal_4340), .Z1_f (new_AGEMA_signal_4341) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4339), .A1_t (new_AGEMA_signal_4340), .A1_f (new_AGEMA_signal_4341), .B0_t (keyFF_outputPar[36]), .B0_f (new_AGEMA_signal_2336), .B1_t (new_AGEMA_signal_2337), .B1_f (new_AGEMA_signal_2338), .Z0_t (keyFF_outputPar[40]), .Z0_f (new_AGEMA_signal_2372), .Z1_t (new_AGEMA_signal_2373), .Z1_f (new_AGEMA_signal_2374) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[37]), .A0_f (new_AGEMA_signal_2345), .A1_t (new_AGEMA_signal_2346), .A1_f (new_AGEMA_signal_2347), .B0_t (keyFF_inputPar[41]), .B0_f (new_AGEMA_signal_3496), .B1_t (new_AGEMA_signal_3497), .B1_f (new_AGEMA_signal_3498), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3905), .Z1_t (new_AGEMA_signal_3906), .Z1_f (new_AGEMA_signal_3907) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3905), .B1_t (new_AGEMA_signal_3906), .B1_f (new_AGEMA_signal_3907), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4342), .Z1_t (new_AGEMA_signal_4343), .Z1_f (new_AGEMA_signal_4344) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4342), .A1_t (new_AGEMA_signal_4343), .A1_f (new_AGEMA_signal_4344), .B0_t (keyFF_outputPar[37]), .B0_f (new_AGEMA_signal_2345), .B1_t (new_AGEMA_signal_2346), .B1_f (new_AGEMA_signal_2347), .Z0_t (keyFF_outputPar[41]), .Z0_f (new_AGEMA_signal_2381), .Z1_t (new_AGEMA_signal_2382), .Z1_f (new_AGEMA_signal_2383) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[38]), .A0_f (new_AGEMA_signal_2354), .A1_t (new_AGEMA_signal_2355), .A1_f (new_AGEMA_signal_2356), .B0_t (keyFF_inputPar[42]), .B0_f (new_AGEMA_signal_3499), .B1_t (new_AGEMA_signal_3500), .B1_f (new_AGEMA_signal_3501), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3908), .Z1_t (new_AGEMA_signal_3909), .Z1_f (new_AGEMA_signal_3910) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3908), .B1_t (new_AGEMA_signal_3909), .B1_f (new_AGEMA_signal_3910), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4345), .Z1_t (new_AGEMA_signal_4346), .Z1_f (new_AGEMA_signal_4347) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4345), .A1_t (new_AGEMA_signal_4346), .A1_f (new_AGEMA_signal_4347), .B0_t (keyFF_outputPar[38]), .B0_f (new_AGEMA_signal_2354), .B1_t (new_AGEMA_signal_2355), .B1_f (new_AGEMA_signal_2356), .Z0_t (keyFF_outputPar[42]), .Z0_f (new_AGEMA_signal_2390), .Z1_t (new_AGEMA_signal_2391), .Z1_f (new_AGEMA_signal_2392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[39]), .A0_f (new_AGEMA_signal_2363), .A1_t (new_AGEMA_signal_2364), .A1_f (new_AGEMA_signal_2365), .B0_t (keyFF_inputPar[43]), .B0_f (new_AGEMA_signal_3502), .B1_t (new_AGEMA_signal_3503), .B1_f (new_AGEMA_signal_3504), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3911), .Z1_t (new_AGEMA_signal_3912), .Z1_f (new_AGEMA_signal_3913) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3911), .B1_t (new_AGEMA_signal_3912), .B1_f (new_AGEMA_signal_3913), .Z0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4348), .Z1_t (new_AGEMA_signal_4349), .Z1_f (new_AGEMA_signal_4350) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4348), .A1_t (new_AGEMA_signal_4349), .A1_f (new_AGEMA_signal_4350), .B0_t (keyFF_outputPar[39]), .B0_f (new_AGEMA_signal_2363), .B1_t (new_AGEMA_signal_2364), .B1_f (new_AGEMA_signal_2365), .Z0_t (keyFF_outputPar[43]), .Z0_f (new_AGEMA_signal_2399), .Z1_t (new_AGEMA_signal_2400), .Z1_f (new_AGEMA_signal_2401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[40]), .A0_f (new_AGEMA_signal_2372), .A1_t (new_AGEMA_signal_2373), .A1_f (new_AGEMA_signal_2374), .B0_t (keyFF_inputPar[44]), .B0_f (new_AGEMA_signal_3505), .B1_t (new_AGEMA_signal_3506), .B1_f (new_AGEMA_signal_3507), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3914), .Z1_t (new_AGEMA_signal_3915), .Z1_f (new_AGEMA_signal_3916) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3914), .B1_t (new_AGEMA_signal_3915), .B1_f (new_AGEMA_signal_3916), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4351), .Z1_t (new_AGEMA_signal_4352), .Z1_f (new_AGEMA_signal_4353) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4351), .A1_t (new_AGEMA_signal_4352), .A1_f (new_AGEMA_signal_4353), .B0_t (keyFF_outputPar[40]), .B0_f (new_AGEMA_signal_2372), .B1_t (new_AGEMA_signal_2373), .B1_f (new_AGEMA_signal_2374), .Z0_t (keyFF_outputPar[44]), .Z0_f (new_AGEMA_signal_2408), .Z1_t (new_AGEMA_signal_2409), .Z1_f (new_AGEMA_signal_2410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[41]), .A0_f (new_AGEMA_signal_2381), .A1_t (new_AGEMA_signal_2382), .A1_f (new_AGEMA_signal_2383), .B0_t (keyFF_inputPar[45]), .B0_f (new_AGEMA_signal_3508), .B1_t (new_AGEMA_signal_3509), .B1_f (new_AGEMA_signal_3510), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3917), .Z1_t (new_AGEMA_signal_3918), .Z1_f (new_AGEMA_signal_3919) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3917), .B1_t (new_AGEMA_signal_3918), .B1_f (new_AGEMA_signal_3919), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4354), .Z1_t (new_AGEMA_signal_4355), .Z1_f (new_AGEMA_signal_4356) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4354), .A1_t (new_AGEMA_signal_4355), .A1_f (new_AGEMA_signal_4356), .B0_t (keyFF_outputPar[41]), .B0_f (new_AGEMA_signal_2381), .B1_t (new_AGEMA_signal_2382), .B1_f (new_AGEMA_signal_2383), .Z0_t (keyFF_outputPar[45]), .Z0_f (new_AGEMA_signal_2417), .Z1_t (new_AGEMA_signal_2418), .Z1_f (new_AGEMA_signal_2419) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[42]), .A0_f (new_AGEMA_signal_2390), .A1_t (new_AGEMA_signal_2391), .A1_f (new_AGEMA_signal_2392), .B0_t (keyFF_inputPar[46]), .B0_f (new_AGEMA_signal_3511), .B1_t (new_AGEMA_signal_3512), .B1_f (new_AGEMA_signal_3513), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3920), .Z1_t (new_AGEMA_signal_3921), .Z1_f (new_AGEMA_signal_3922) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3920), .B1_t (new_AGEMA_signal_3921), .B1_f (new_AGEMA_signal_3922), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4357), .Z1_t (new_AGEMA_signal_4358), .Z1_f (new_AGEMA_signal_4359) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4357), .A1_t (new_AGEMA_signal_4358), .A1_f (new_AGEMA_signal_4359), .B0_t (keyFF_outputPar[42]), .B0_f (new_AGEMA_signal_2390), .B1_t (new_AGEMA_signal_2391), .B1_f (new_AGEMA_signal_2392), .Z0_t (keyFF_outputPar[46]), .Z0_f (new_AGEMA_signal_2426), .Z1_t (new_AGEMA_signal_2427), .Z1_f (new_AGEMA_signal_2428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[43]), .A0_f (new_AGEMA_signal_2399), .A1_t (new_AGEMA_signal_2400), .A1_f (new_AGEMA_signal_2401), .B0_t (keyFF_inputPar[47]), .B0_f (new_AGEMA_signal_3514), .B1_t (new_AGEMA_signal_3515), .B1_f (new_AGEMA_signal_3516), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3923), .Z1_t (new_AGEMA_signal_3924), .Z1_f (new_AGEMA_signal_3925) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3923), .B1_t (new_AGEMA_signal_3924), .B1_f (new_AGEMA_signal_3925), .Z0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4360), .Z1_t (new_AGEMA_signal_4361), .Z1_f (new_AGEMA_signal_4362) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4360), .A1_t (new_AGEMA_signal_4361), .A1_f (new_AGEMA_signal_4362), .B0_t (keyFF_outputPar[43]), .B0_f (new_AGEMA_signal_2399), .B1_t (new_AGEMA_signal_2400), .B1_f (new_AGEMA_signal_2401), .Z0_t (keyFF_outputPar[47]), .Z0_f (new_AGEMA_signal_2435), .Z1_t (new_AGEMA_signal_2436), .Z1_f (new_AGEMA_signal_2437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[44]), .A0_f (new_AGEMA_signal_2408), .A1_t (new_AGEMA_signal_2409), .A1_f (new_AGEMA_signal_2410), .B0_t (keyFF_inputPar[48]), .B0_f (new_AGEMA_signal_3517), .B1_t (new_AGEMA_signal_3518), .B1_f (new_AGEMA_signal_3519), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3926), .Z1_t (new_AGEMA_signal_3927), .Z1_f (new_AGEMA_signal_3928) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3926), .B1_t (new_AGEMA_signal_3927), .B1_f (new_AGEMA_signal_3928), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4363), .Z1_t (new_AGEMA_signal_4364), .Z1_f (new_AGEMA_signal_4365) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4363), .A1_t (new_AGEMA_signal_4364), .A1_f (new_AGEMA_signal_4365), .B0_t (keyFF_outputPar[44]), .B0_f (new_AGEMA_signal_2408), .B1_t (new_AGEMA_signal_2409), .B1_f (new_AGEMA_signal_2410), .Z0_t (keyFF_outputPar[48]), .Z0_f (new_AGEMA_signal_2444), .Z1_t (new_AGEMA_signal_2445), .Z1_f (new_AGEMA_signal_2446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[45]), .A0_f (new_AGEMA_signal_2417), .A1_t (new_AGEMA_signal_2418), .A1_f (new_AGEMA_signal_2419), .B0_t (keyFF_inputPar[49]), .B0_f (new_AGEMA_signal_3520), .B1_t (new_AGEMA_signal_3521), .B1_f (new_AGEMA_signal_3522), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3929), .Z1_t (new_AGEMA_signal_3930), .Z1_f (new_AGEMA_signal_3931) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3929), .B1_t (new_AGEMA_signal_3930), .B1_f (new_AGEMA_signal_3931), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4366), .Z1_t (new_AGEMA_signal_4367), .Z1_f (new_AGEMA_signal_4368) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4366), .A1_t (new_AGEMA_signal_4367), .A1_f (new_AGEMA_signal_4368), .B0_t (keyFF_outputPar[45]), .B0_f (new_AGEMA_signal_2417), .B1_t (new_AGEMA_signal_2418), .B1_f (new_AGEMA_signal_2419), .Z0_t (keyFF_outputPar[49]), .Z0_f (new_AGEMA_signal_2453), .Z1_t (new_AGEMA_signal_2454), .Z1_f (new_AGEMA_signal_2455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[46]), .A0_f (new_AGEMA_signal_2426), .A1_t (new_AGEMA_signal_2427), .A1_f (new_AGEMA_signal_2428), .B0_t (keyFF_inputPar[50]), .B0_f (new_AGEMA_signal_3523), .B1_t (new_AGEMA_signal_3524), .B1_f (new_AGEMA_signal_3525), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3932), .Z1_t (new_AGEMA_signal_3933), .Z1_f (new_AGEMA_signal_3934) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3932), .B1_t (new_AGEMA_signal_3933), .B1_f (new_AGEMA_signal_3934), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4369), .Z1_t (new_AGEMA_signal_4370), .Z1_f (new_AGEMA_signal_4371) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4369), .A1_t (new_AGEMA_signal_4370), .A1_f (new_AGEMA_signal_4371), .B0_t (keyFF_outputPar[46]), .B0_f (new_AGEMA_signal_2426), .B1_t (new_AGEMA_signal_2427), .B1_f (new_AGEMA_signal_2428), .Z0_t (keyFF_outputPar[50]), .Z0_f (new_AGEMA_signal_2462), .Z1_t (new_AGEMA_signal_2463), .Z1_f (new_AGEMA_signal_2464) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[47]), .A0_f (new_AGEMA_signal_2435), .A1_t (new_AGEMA_signal_2436), .A1_f (new_AGEMA_signal_2437), .B0_t (keyFF_inputPar[51]), .B0_f (new_AGEMA_signal_3526), .B1_t (new_AGEMA_signal_3527), .B1_f (new_AGEMA_signal_3528), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3935), .Z1_t (new_AGEMA_signal_3936), .Z1_f (new_AGEMA_signal_3937) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3935), .B1_t (new_AGEMA_signal_3936), .B1_f (new_AGEMA_signal_3937), .Z0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4372), .Z1_t (new_AGEMA_signal_4373), .Z1_f (new_AGEMA_signal_4374) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4372), .A1_t (new_AGEMA_signal_4373), .A1_f (new_AGEMA_signal_4374), .B0_t (keyFF_outputPar[47]), .B0_f (new_AGEMA_signal_2435), .B1_t (new_AGEMA_signal_2436), .B1_f (new_AGEMA_signal_2437), .Z0_t (keyFF_outputPar[51]), .Z0_f (new_AGEMA_signal_2471), .Z1_t (new_AGEMA_signal_2472), .Z1_f (new_AGEMA_signal_2473) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[48]), .A0_f (new_AGEMA_signal_2444), .A1_t (new_AGEMA_signal_2445), .A1_f (new_AGEMA_signal_2446), .B0_t (keyFF_inputPar[52]), .B0_f (new_AGEMA_signal_3529), .B1_t (new_AGEMA_signal_3530), .B1_f (new_AGEMA_signal_3531), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3938), .Z1_t (new_AGEMA_signal_3939), .Z1_f (new_AGEMA_signal_3940) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3938), .B1_t (new_AGEMA_signal_3939), .B1_f (new_AGEMA_signal_3940), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4375), .Z1_t (new_AGEMA_signal_4376), .Z1_f (new_AGEMA_signal_4377) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4375), .A1_t (new_AGEMA_signal_4376), .A1_f (new_AGEMA_signal_4377), .B0_t (keyFF_outputPar[48]), .B0_f (new_AGEMA_signal_2444), .B1_t (new_AGEMA_signal_2445), .B1_f (new_AGEMA_signal_2446), .Z0_t (keyFF_outputPar[52]), .Z0_f (new_AGEMA_signal_2480), .Z1_t (new_AGEMA_signal_2481), .Z1_f (new_AGEMA_signal_2482) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[49]), .A0_f (new_AGEMA_signal_2453), .A1_t (new_AGEMA_signal_2454), .A1_f (new_AGEMA_signal_2455), .B0_t (keyFF_inputPar[53]), .B0_f (new_AGEMA_signal_3532), .B1_t (new_AGEMA_signal_3533), .B1_f (new_AGEMA_signal_3534), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3941), .Z1_t (new_AGEMA_signal_3942), .Z1_f (new_AGEMA_signal_3943) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3941), .B1_t (new_AGEMA_signal_3942), .B1_f (new_AGEMA_signal_3943), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4378), .Z1_t (new_AGEMA_signal_4379), .Z1_f (new_AGEMA_signal_4380) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4378), .A1_t (new_AGEMA_signal_4379), .A1_f (new_AGEMA_signal_4380), .B0_t (keyFF_outputPar[49]), .B0_f (new_AGEMA_signal_2453), .B1_t (new_AGEMA_signal_2454), .B1_f (new_AGEMA_signal_2455), .Z0_t (keyFF_outputPar[53]), .Z0_f (new_AGEMA_signal_2489), .Z1_t (new_AGEMA_signal_2490), .Z1_f (new_AGEMA_signal_2491) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[50]), .A0_f (new_AGEMA_signal_2462), .A1_t (new_AGEMA_signal_2463), .A1_f (new_AGEMA_signal_2464), .B0_t (keyFF_inputPar[54]), .B0_f (new_AGEMA_signal_3535), .B1_t (new_AGEMA_signal_3536), .B1_f (new_AGEMA_signal_3537), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3944), .Z1_t (new_AGEMA_signal_3945), .Z1_f (new_AGEMA_signal_3946) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3944), .B1_t (new_AGEMA_signal_3945), .B1_f (new_AGEMA_signal_3946), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4381), .Z1_t (new_AGEMA_signal_4382), .Z1_f (new_AGEMA_signal_4383) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4381), .A1_t (new_AGEMA_signal_4382), .A1_f (new_AGEMA_signal_4383), .B0_t (keyFF_outputPar[50]), .B0_f (new_AGEMA_signal_2462), .B1_t (new_AGEMA_signal_2463), .B1_f (new_AGEMA_signal_2464), .Z0_t (keyFF_outputPar[54]), .Z0_f (new_AGEMA_signal_2498), .Z1_t (new_AGEMA_signal_2499), .Z1_f (new_AGEMA_signal_2500) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[51]), .A0_f (new_AGEMA_signal_2471), .A1_t (new_AGEMA_signal_2472), .A1_f (new_AGEMA_signal_2473), .B0_t (keyFF_inputPar[55]), .B0_f (new_AGEMA_signal_3538), .B1_t (new_AGEMA_signal_3539), .B1_f (new_AGEMA_signal_3540), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3947), .Z1_t (new_AGEMA_signal_3948), .Z1_f (new_AGEMA_signal_3949) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3947), .B1_t (new_AGEMA_signal_3948), .B1_f (new_AGEMA_signal_3949), .Z0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4384), .Z1_t (new_AGEMA_signal_4385), .Z1_f (new_AGEMA_signal_4386) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4384), .A1_t (new_AGEMA_signal_4385), .A1_f (new_AGEMA_signal_4386), .B0_t (keyFF_outputPar[51]), .B0_f (new_AGEMA_signal_2471), .B1_t (new_AGEMA_signal_2472), .B1_f (new_AGEMA_signal_2473), .Z0_t (keyFF_outputPar[55]), .Z0_f (new_AGEMA_signal_2507), .Z1_t (new_AGEMA_signal_2508), .Z1_f (new_AGEMA_signal_2509) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[52]), .A0_f (new_AGEMA_signal_2480), .A1_t (new_AGEMA_signal_2481), .A1_f (new_AGEMA_signal_2482), .B0_t (keyFF_inputPar[56]), .B0_f (new_AGEMA_signal_3541), .B1_t (new_AGEMA_signal_3542), .B1_f (new_AGEMA_signal_3543), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3950), .Z1_t (new_AGEMA_signal_3951), .Z1_f (new_AGEMA_signal_3952) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3950), .B1_t (new_AGEMA_signal_3951), .B1_f (new_AGEMA_signal_3952), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4387), .Z1_t (new_AGEMA_signal_4388), .Z1_f (new_AGEMA_signal_4389) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4387), .A1_t (new_AGEMA_signal_4388), .A1_f (new_AGEMA_signal_4389), .B0_t (keyFF_outputPar[52]), .B0_f (new_AGEMA_signal_2480), .B1_t (new_AGEMA_signal_2481), .B1_f (new_AGEMA_signal_2482), .Z0_t (keyFF_outputPar[56]), .Z0_f (new_AGEMA_signal_2516), .Z1_t (new_AGEMA_signal_2517), .Z1_f (new_AGEMA_signal_2518) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[53]), .A0_f (new_AGEMA_signal_2489), .A1_t (new_AGEMA_signal_2490), .A1_f (new_AGEMA_signal_2491), .B0_t (keyFF_inputPar[57]), .B0_f (new_AGEMA_signal_3544), .B1_t (new_AGEMA_signal_3545), .B1_f (new_AGEMA_signal_3546), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3953), .Z1_t (new_AGEMA_signal_3954), .Z1_f (new_AGEMA_signal_3955) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3953), .B1_t (new_AGEMA_signal_3954), .B1_f (new_AGEMA_signal_3955), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4390), .Z1_t (new_AGEMA_signal_4391), .Z1_f (new_AGEMA_signal_4392) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4390), .A1_t (new_AGEMA_signal_4391), .A1_f (new_AGEMA_signal_4392), .B0_t (keyFF_outputPar[53]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (keyFF_outputPar[57]), .Z0_f (new_AGEMA_signal_2525), .Z1_t (new_AGEMA_signal_2526), .Z1_f (new_AGEMA_signal_2527) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[54]), .A0_f (new_AGEMA_signal_2498), .A1_t (new_AGEMA_signal_2499), .A1_f (new_AGEMA_signal_2500), .B0_t (keyFF_inputPar[58]), .B0_f (new_AGEMA_signal_3547), .B1_t (new_AGEMA_signal_3548), .B1_f (new_AGEMA_signal_3549), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3956), .Z1_t (new_AGEMA_signal_3957), .Z1_f (new_AGEMA_signal_3958) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3956), .B1_t (new_AGEMA_signal_3957), .B1_f (new_AGEMA_signal_3958), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4393), .Z1_t (new_AGEMA_signal_4394), .Z1_f (new_AGEMA_signal_4395) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4393), .A1_t (new_AGEMA_signal_4394), .A1_f (new_AGEMA_signal_4395), .B0_t (keyFF_outputPar[54]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (keyFF_outputPar[58]), .Z0_f (new_AGEMA_signal_2534), .Z1_t (new_AGEMA_signal_2535), .Z1_f (new_AGEMA_signal_2536) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[55]), .A0_f (new_AGEMA_signal_2507), .A1_t (new_AGEMA_signal_2508), .A1_f (new_AGEMA_signal_2509), .B0_t (keyFF_inputPar[59]), .B0_f (new_AGEMA_signal_3550), .B1_t (new_AGEMA_signal_3551), .B1_f (new_AGEMA_signal_3552), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3959), .Z1_t (new_AGEMA_signal_3960), .Z1_f (new_AGEMA_signal_3961) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3959), .B1_t (new_AGEMA_signal_3960), .B1_f (new_AGEMA_signal_3961), .Z0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4396), .Z1_t (new_AGEMA_signal_4397), .Z1_f (new_AGEMA_signal_4398) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4396), .A1_t (new_AGEMA_signal_4397), .A1_f (new_AGEMA_signal_4398), .B0_t (keyFF_outputPar[55]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (keyFF_outputPar[59]), .Z0_f (new_AGEMA_signal_2543), .Z1_t (new_AGEMA_signal_2544), .Z1_f (new_AGEMA_signal_2545) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[56]), .A0_f (new_AGEMA_signal_2516), .A1_t (new_AGEMA_signal_2517), .A1_f (new_AGEMA_signal_2518), .B0_t (keyFF_inputPar[60]), .B0_f (new_AGEMA_signal_3553), .B1_t (new_AGEMA_signal_3554), .B1_f (new_AGEMA_signal_3555), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3962), .Z1_t (new_AGEMA_signal_3963), .Z1_f (new_AGEMA_signal_3964) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3962), .B1_t (new_AGEMA_signal_3963), .B1_f (new_AGEMA_signal_3964), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4399), .Z1_t (new_AGEMA_signal_4400), .Z1_f (new_AGEMA_signal_4401) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4399), .A1_t (new_AGEMA_signal_4400), .A1_f (new_AGEMA_signal_4401), .B0_t (keyFF_outputPar[56]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (keyFF_outputPar[60]), .Z0_f (new_AGEMA_signal_2552), .Z1_t (new_AGEMA_signal_2553), .Z1_f (new_AGEMA_signal_2554) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[57]), .A0_f (new_AGEMA_signal_2525), .A1_t (new_AGEMA_signal_2526), .A1_f (new_AGEMA_signal_2527), .B0_t (keyFF_inputPar[61]), .B0_f (new_AGEMA_signal_3556), .B1_t (new_AGEMA_signal_3557), .B1_f (new_AGEMA_signal_3558), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3965), .Z1_t (new_AGEMA_signal_3966), .Z1_f (new_AGEMA_signal_3967) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3965), .B1_t (new_AGEMA_signal_3966), .B1_f (new_AGEMA_signal_3967), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4402), .Z1_t (new_AGEMA_signal_4403), .Z1_f (new_AGEMA_signal_4404) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4402), .A1_t (new_AGEMA_signal_4403), .A1_f (new_AGEMA_signal_4404), .B0_t (keyFF_outputPar[57]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (keyFF_outputPar[61]), .Z0_f (new_AGEMA_signal_2561), .Z1_t (new_AGEMA_signal_2562), .Z1_f (new_AGEMA_signal_2563) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[58]), .A0_f (new_AGEMA_signal_2534), .A1_t (new_AGEMA_signal_2535), .A1_f (new_AGEMA_signal_2536), .B0_t (keyFF_inputPar[62]), .B0_f (new_AGEMA_signal_3559), .B1_t (new_AGEMA_signal_3560), .B1_f (new_AGEMA_signal_3561), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3968), .Z1_t (new_AGEMA_signal_3969), .Z1_f (new_AGEMA_signal_3970) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3968), .B1_t (new_AGEMA_signal_3969), .B1_f (new_AGEMA_signal_3970), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4405), .Z1_t (new_AGEMA_signal_4406), .Z1_f (new_AGEMA_signal_4407) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4405), .A1_t (new_AGEMA_signal_4406), .A1_f (new_AGEMA_signal_4407), .B0_t (keyFF_outputPar[58]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (keyFF_outputPar[62]), .Z0_f (new_AGEMA_signal_2570), .Z1_t (new_AGEMA_signal_2571), .Z1_f (new_AGEMA_signal_2572) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[59]), .A0_f (new_AGEMA_signal_2543), .A1_t (new_AGEMA_signal_2544), .A1_f (new_AGEMA_signal_2545), .B0_t (keyFF_inputPar[63]), .B0_f (new_AGEMA_signal_3562), .B1_t (new_AGEMA_signal_3563), .B1_f (new_AGEMA_signal_3564), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3971), .Z1_t (new_AGEMA_signal_3972), .Z1_f (new_AGEMA_signal_3973) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3971), .B1_t (new_AGEMA_signal_3972), .B1_f (new_AGEMA_signal_3973), .Z0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4408), .Z1_t (new_AGEMA_signal_4409), .Z1_f (new_AGEMA_signal_4410) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4408), .A1_t (new_AGEMA_signal_4409), .A1_f (new_AGEMA_signal_4410), .B0_t (keyFF_outputPar[59]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (keyFF_outputPar[63]), .Z0_f (new_AGEMA_signal_2579), .Z1_t (new_AGEMA_signal_2580), .Z1_f (new_AGEMA_signal_2581) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[60]), .A0_f (new_AGEMA_signal_2552), .A1_t (new_AGEMA_signal_2553), .A1_f (new_AGEMA_signal_2554), .B0_t (keyFF_inputPar[64]), .B0_f (new_AGEMA_signal_3565), .B1_t (new_AGEMA_signal_3566), .B1_f (new_AGEMA_signal_3567), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3974), .Z1_t (new_AGEMA_signal_3975), .Z1_f (new_AGEMA_signal_3976) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3974), .B1_t (new_AGEMA_signal_3975), .B1_f (new_AGEMA_signal_3976), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4411), .Z1_t (new_AGEMA_signal_4412), .Z1_f (new_AGEMA_signal_4413) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4411), .A1_t (new_AGEMA_signal_4412), .A1_f (new_AGEMA_signal_4413), .B0_t (keyFF_outputPar[60]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (keyFF_outputPar[64]), .Z0_f (new_AGEMA_signal_2588), .Z1_t (new_AGEMA_signal_2589), .Z1_f (new_AGEMA_signal_2590) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[61]), .A0_f (new_AGEMA_signal_2561), .A1_t (new_AGEMA_signal_2562), .A1_f (new_AGEMA_signal_2563), .B0_t (keyFF_inputPar[65]), .B0_f (new_AGEMA_signal_3568), .B1_t (new_AGEMA_signal_3569), .B1_f (new_AGEMA_signal_3570), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3977), .Z1_t (new_AGEMA_signal_3978), .Z1_f (new_AGEMA_signal_3979) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3977), .B1_t (new_AGEMA_signal_3978), .B1_f (new_AGEMA_signal_3979), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4414), .Z1_t (new_AGEMA_signal_4415), .Z1_f (new_AGEMA_signal_4416) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4414), .A1_t (new_AGEMA_signal_4415), .A1_f (new_AGEMA_signal_4416), .B0_t (keyFF_outputPar[61]), .B0_f (new_AGEMA_signal_2561), .B1_t (new_AGEMA_signal_2562), .B1_f (new_AGEMA_signal_2563), .Z0_t (keyFF_outputPar[65]), .Z0_f (new_AGEMA_signal_2597), .Z1_t (new_AGEMA_signal_2598), .Z1_f (new_AGEMA_signal_2599) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[62]), .A0_f (new_AGEMA_signal_2570), .A1_t (new_AGEMA_signal_2571), .A1_f (new_AGEMA_signal_2572), .B0_t (keyFF_inputPar[66]), .B0_f (new_AGEMA_signal_3571), .B1_t (new_AGEMA_signal_3572), .B1_f (new_AGEMA_signal_3573), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3980), .Z1_t (new_AGEMA_signal_3981), .Z1_f (new_AGEMA_signal_3982) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3980), .B1_t (new_AGEMA_signal_3981), .B1_f (new_AGEMA_signal_3982), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4417), .Z1_t (new_AGEMA_signal_4418), .Z1_f (new_AGEMA_signal_4419) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4417), .A1_t (new_AGEMA_signal_4418), .A1_f (new_AGEMA_signal_4419), .B0_t (keyFF_outputPar[62]), .B0_f (new_AGEMA_signal_2570), .B1_t (new_AGEMA_signal_2571), .B1_f (new_AGEMA_signal_2572), .Z0_t (keyFF_outputPar[66]), .Z0_f (new_AGEMA_signal_2606), .Z1_t (new_AGEMA_signal_2607), .Z1_f (new_AGEMA_signal_2608) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[63]), .A0_f (new_AGEMA_signal_2579), .A1_t (new_AGEMA_signal_2580), .A1_f (new_AGEMA_signal_2581), .B0_t (keyFF_inputPar[67]), .B0_f (new_AGEMA_signal_3574), .B1_t (new_AGEMA_signal_3575), .B1_f (new_AGEMA_signal_3576), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3983), .Z1_t (new_AGEMA_signal_3984), .Z1_f (new_AGEMA_signal_3985) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3983), .B1_t (new_AGEMA_signal_3984), .B1_f (new_AGEMA_signal_3985), .Z0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4420), .Z1_t (new_AGEMA_signal_4421), .Z1_f (new_AGEMA_signal_4422) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4420), .A1_t (new_AGEMA_signal_4421), .A1_f (new_AGEMA_signal_4422), .B0_t (keyFF_outputPar[63]), .B0_f (new_AGEMA_signal_2579), .B1_t (new_AGEMA_signal_2580), .B1_f (new_AGEMA_signal_2581), .Z0_t (keyFF_outputPar[67]), .Z0_f (new_AGEMA_signal_2615), .Z1_t (new_AGEMA_signal_2616), .Z1_f (new_AGEMA_signal_2617) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[64]), .A0_f (new_AGEMA_signal_2588), .A1_t (new_AGEMA_signal_2589), .A1_f (new_AGEMA_signal_2590), .B0_t (keyFF_inputPar[68]), .B0_f (new_AGEMA_signal_3577), .B1_t (new_AGEMA_signal_3578), .B1_f (new_AGEMA_signal_3579), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3986), .Z1_t (new_AGEMA_signal_3987), .Z1_f (new_AGEMA_signal_3988) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3986), .B1_t (new_AGEMA_signal_3987), .B1_f (new_AGEMA_signal_3988), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4423), .Z1_t (new_AGEMA_signal_4424), .Z1_f (new_AGEMA_signal_4425) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4423), .A1_t (new_AGEMA_signal_4424), .A1_f (new_AGEMA_signal_4425), .B0_t (keyFF_outputPar[64]), .B0_f (new_AGEMA_signal_2588), .B1_t (new_AGEMA_signal_2589), .B1_f (new_AGEMA_signal_2590), .Z0_t (keyFF_outputPar[68]), .Z0_f (new_AGEMA_signal_2624), .Z1_t (new_AGEMA_signal_2625), .Z1_f (new_AGEMA_signal_2626) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[65]), .A0_f (new_AGEMA_signal_2597), .A1_t (new_AGEMA_signal_2598), .A1_f (new_AGEMA_signal_2599), .B0_t (keyFF_inputPar[69]), .B0_f (new_AGEMA_signal_3580), .B1_t (new_AGEMA_signal_3581), .B1_f (new_AGEMA_signal_3582), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3989), .Z1_t (new_AGEMA_signal_3990), .Z1_f (new_AGEMA_signal_3991) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3989), .B1_t (new_AGEMA_signal_3990), .B1_f (new_AGEMA_signal_3991), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4426), .Z1_t (new_AGEMA_signal_4427), .Z1_f (new_AGEMA_signal_4428) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4426), .A1_t (new_AGEMA_signal_4427), .A1_f (new_AGEMA_signal_4428), .B0_t (keyFF_outputPar[65]), .B0_f (new_AGEMA_signal_2597), .B1_t (new_AGEMA_signal_2598), .B1_f (new_AGEMA_signal_2599), .Z0_t (keyFF_outputPar[69]), .Z0_f (new_AGEMA_signal_2633), .Z1_t (new_AGEMA_signal_2634), .Z1_f (new_AGEMA_signal_2635) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[66]), .A0_f (new_AGEMA_signal_2606), .A1_t (new_AGEMA_signal_2607), .A1_f (new_AGEMA_signal_2608), .B0_t (keyFF_inputPar[70]), .B0_f (new_AGEMA_signal_3583), .B1_t (new_AGEMA_signal_3584), .B1_f (new_AGEMA_signal_3585), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3992), .Z1_t (new_AGEMA_signal_3993), .Z1_f (new_AGEMA_signal_3994) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3992), .B1_t (new_AGEMA_signal_3993), .B1_f (new_AGEMA_signal_3994), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4429), .Z1_t (new_AGEMA_signal_4430), .Z1_f (new_AGEMA_signal_4431) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4429), .A1_t (new_AGEMA_signal_4430), .A1_f (new_AGEMA_signal_4431), .B0_t (keyFF_outputPar[66]), .B0_f (new_AGEMA_signal_2606), .B1_t (new_AGEMA_signal_2607), .B1_f (new_AGEMA_signal_2608), .Z0_t (keyFF_outputPar[70]), .Z0_f (new_AGEMA_signal_2642), .Z1_t (new_AGEMA_signal_2643), .Z1_f (new_AGEMA_signal_2644) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[67]), .A0_f (new_AGEMA_signal_2615), .A1_t (new_AGEMA_signal_2616), .A1_f (new_AGEMA_signal_2617), .B0_t (keyFF_inputPar[71]), .B0_f (new_AGEMA_signal_3586), .B1_t (new_AGEMA_signal_3587), .B1_f (new_AGEMA_signal_3588), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3995), .Z1_t (new_AGEMA_signal_3996), .Z1_f (new_AGEMA_signal_3997) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3995), .B1_t (new_AGEMA_signal_3996), .B1_f (new_AGEMA_signal_3997), .Z0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4432), .Z1_t (new_AGEMA_signal_4433), .Z1_f (new_AGEMA_signal_4434) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4432), .A1_t (new_AGEMA_signal_4433), .A1_f (new_AGEMA_signal_4434), .B0_t (keyFF_outputPar[67]), .B0_f (new_AGEMA_signal_2615), .B1_t (new_AGEMA_signal_2616), .B1_f (new_AGEMA_signal_2617), .Z0_t (keyFF_outputPar[71]), .Z0_f (new_AGEMA_signal_2651), .Z1_t (new_AGEMA_signal_2652), .Z1_f (new_AGEMA_signal_2653) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[68]), .A0_f (new_AGEMA_signal_2624), .A1_t (new_AGEMA_signal_2625), .A1_f (new_AGEMA_signal_2626), .B0_t (keyFF_inputPar[72]), .B0_f (new_AGEMA_signal_3589), .B1_t (new_AGEMA_signal_3590), .B1_f (new_AGEMA_signal_3591), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3998), .Z1_t (new_AGEMA_signal_3999), .Z1_f (new_AGEMA_signal_4000) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3998), .B1_t (new_AGEMA_signal_3999), .B1_f (new_AGEMA_signal_4000), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4435), .Z1_t (new_AGEMA_signal_4436), .Z1_f (new_AGEMA_signal_4437) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4435), .A1_t (new_AGEMA_signal_4436), .A1_f (new_AGEMA_signal_4437), .B0_t (keyFF_outputPar[68]), .B0_f (new_AGEMA_signal_2624), .B1_t (new_AGEMA_signal_2625), .B1_f (new_AGEMA_signal_2626), .Z0_t (keyFF_outputPar[72]), .Z0_f (new_AGEMA_signal_2660), .Z1_t (new_AGEMA_signal_2661), .Z1_f (new_AGEMA_signal_2662) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[69]), .A0_f (new_AGEMA_signal_2633), .A1_t (new_AGEMA_signal_2634), .A1_f (new_AGEMA_signal_2635), .B0_t (keyFF_inputPar[73]), .B0_f (new_AGEMA_signal_3592), .B1_t (new_AGEMA_signal_3593), .B1_f (new_AGEMA_signal_3594), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4001), .Z1_t (new_AGEMA_signal_4002), .Z1_f (new_AGEMA_signal_4003) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4001), .B1_t (new_AGEMA_signal_4002), .B1_f (new_AGEMA_signal_4003), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4438), .Z1_t (new_AGEMA_signal_4439), .Z1_f (new_AGEMA_signal_4440) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4438), .A1_t (new_AGEMA_signal_4439), .A1_f (new_AGEMA_signal_4440), .B0_t (keyFF_outputPar[69]), .B0_f (new_AGEMA_signal_2633), .B1_t (new_AGEMA_signal_2634), .B1_f (new_AGEMA_signal_2635), .Z0_t (keyFF_outputPar[73]), .Z0_f (new_AGEMA_signal_2669), .Z1_t (new_AGEMA_signal_2670), .Z1_f (new_AGEMA_signal_2671) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[70]), .A0_f (new_AGEMA_signal_2642), .A1_t (new_AGEMA_signal_2643), .A1_f (new_AGEMA_signal_2644), .B0_t (keyFF_inputPar[74]), .B0_f (new_AGEMA_signal_3595), .B1_t (new_AGEMA_signal_3596), .B1_f (new_AGEMA_signal_3597), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_4004), .Z1_t (new_AGEMA_signal_4005), .Z1_f (new_AGEMA_signal_4006) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_4004), .B1_t (new_AGEMA_signal_4005), .B1_f (new_AGEMA_signal_4006), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4441), .Z1_t (new_AGEMA_signal_4442), .Z1_f (new_AGEMA_signal_4443) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4441), .A1_t (new_AGEMA_signal_4442), .A1_f (new_AGEMA_signal_4443), .B0_t (keyFF_outputPar[70]), .B0_f (new_AGEMA_signal_2642), .B1_t (new_AGEMA_signal_2643), .B1_f (new_AGEMA_signal_2644), .Z0_t (keyFF_outputPar[74]), .Z0_f (new_AGEMA_signal_2678), .Z1_t (new_AGEMA_signal_2679), .Z1_f (new_AGEMA_signal_2680) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[71]), .A0_f (new_AGEMA_signal_2651), .A1_t (new_AGEMA_signal_2652), .A1_f (new_AGEMA_signal_2653), .B0_t (keyFF_inputPar[75]), .B0_f (new_AGEMA_signal_3598), .B1_t (new_AGEMA_signal_3599), .B1_f (new_AGEMA_signal_3600), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4007), .Z1_t (new_AGEMA_signal_4008), .Z1_f (new_AGEMA_signal_4009) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4007), .B1_t (new_AGEMA_signal_4008), .B1_f (new_AGEMA_signal_4009), .Z0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4444), .Z1_t (new_AGEMA_signal_4445), .Z1_f (new_AGEMA_signal_4446) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4444), .A1_t (new_AGEMA_signal_4445), .A1_f (new_AGEMA_signal_4446), .B0_t (keyFF_outputPar[71]), .B0_f (new_AGEMA_signal_2651), .B1_t (new_AGEMA_signal_2652), .B1_f (new_AGEMA_signal_2653), .Z0_t (keyFF_outputPar[75]), .Z0_f (new_AGEMA_signal_2687), .Z1_t (new_AGEMA_signal_2688), .Z1_f (new_AGEMA_signal_2689) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[72]), .A0_f (new_AGEMA_signal_2660), .A1_t (new_AGEMA_signal_2661), .A1_f (new_AGEMA_signal_2662), .B0_t (keyFF_inputPar[76]), .B0_f (new_AGEMA_signal_4526), .B1_t (new_AGEMA_signal_4527), .B1_f (new_AGEMA_signal_4528), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_4541), .Z1_t (new_AGEMA_signal_4542), .Z1_f (new_AGEMA_signal_4543) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_4541), .B1_t (new_AGEMA_signal_4542), .B1_f (new_AGEMA_signal_4543), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4556), .Z1_t (new_AGEMA_signal_4557), .Z1_f (new_AGEMA_signal_4558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4556), .A1_t (new_AGEMA_signal_4557), .A1_f (new_AGEMA_signal_4558), .B0_t (keyFF_outputPar[72]), .B0_f (new_AGEMA_signal_2660), .B1_t (new_AGEMA_signal_2661), .B1_f (new_AGEMA_signal_2662), .Z0_t (roundkey[0]), .Z0_f (new_AGEMA_signal_1452), .Z1_t (new_AGEMA_signal_1453), .Z1_f (new_AGEMA_signal_1454) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[73]), .A0_f (new_AGEMA_signal_2669), .A1_t (new_AGEMA_signal_2670), .A1_f (new_AGEMA_signal_2671), .B0_t (keyFF_inputPar[77]), .B0_f (new_AGEMA_signal_4601), .B1_t (new_AGEMA_signal_4602), .B1_f (new_AGEMA_signal_4603), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4625), .Z1_t (new_AGEMA_signal_4626), .Z1_f (new_AGEMA_signal_4627) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4625), .B1_t (new_AGEMA_signal_4626), .B1_f (new_AGEMA_signal_4627), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4646), .Z1_t (new_AGEMA_signal_4647), .Z1_f (new_AGEMA_signal_4648) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4646), .A1_t (new_AGEMA_signal_4647), .A1_f (new_AGEMA_signal_4648), .B0_t (keyFF_outputPar[73]), .B0_f (new_AGEMA_signal_2669), .B1_t (new_AGEMA_signal_2670), .B1_f (new_AGEMA_signal_2671), .Z0_t (roundkey[1]), .Z0_f (new_AGEMA_signal_1434), .Z1_t (new_AGEMA_signal_1435), .Z1_f (new_AGEMA_signal_1436) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[74]), .A0_f (new_AGEMA_signal_2678), .A1_t (new_AGEMA_signal_2679), .A1_f (new_AGEMA_signal_2680), .B0_t (keyFF_inputPar[78]), .B0_f (new_AGEMA_signal_4604), .B1_t (new_AGEMA_signal_4605), .B1_f (new_AGEMA_signal_4606), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_4628), .Z1_t (new_AGEMA_signal_4629), .Z1_f (new_AGEMA_signal_4630) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_4628), .B1_t (new_AGEMA_signal_4629), .B1_f (new_AGEMA_signal_4630), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4649), .Z1_t (new_AGEMA_signal_4650), .Z1_f (new_AGEMA_signal_4651) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4649), .A1_t (new_AGEMA_signal_4650), .A1_f (new_AGEMA_signal_4651), .B0_t (keyFF_outputPar[74]), .B0_f (new_AGEMA_signal_2678), .B1_t (new_AGEMA_signal_2679), .B1_f (new_AGEMA_signal_2680), .Z0_t (roundkey[2]), .Z0_f (new_AGEMA_signal_1443), .Z1_t (new_AGEMA_signal_1444), .Z1_f (new_AGEMA_signal_1445) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[75]), .A0_f (new_AGEMA_signal_2687), .A1_t (new_AGEMA_signal_2688), .A1_f (new_AGEMA_signal_2689), .B0_t (keyFF_inputPar[79]), .B0_f (new_AGEMA_signal_4631), .B1_t (new_AGEMA_signal_4632), .B1_f (new_AGEMA_signal_4633), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4652), .Z1_t (new_AGEMA_signal_4653), .Z1_f (new_AGEMA_signal_4654) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (fsm_rst_countSerial), .A1_f (new_AGEMA_signal_2717), .B0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4652), .B1_t (new_AGEMA_signal_4653), .B1_f (new_AGEMA_signal_4654), .Z0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4658), .Z1_t (new_AGEMA_signal_4659), .Z1_f (new_AGEMA_signal_4660) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4658), .A1_t (new_AGEMA_signal_4659), .A1_f (new_AGEMA_signal_4660), .B0_t (keyFF_outputPar[75]), .B0_f (new_AGEMA_signal_2687), .B1_t (new_AGEMA_signal_2688), .B1_f (new_AGEMA_signal_2689), .Z0_t (roundkey[3]), .Z0_f (new_AGEMA_signal_1461), .Z1_t (new_AGEMA_signal_1462), .Z1_f (new_AGEMA_signal_1463) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[3]), .A0_f (new_AGEMA_signal_2084), .A1_t (new_AGEMA_signal_2085), .A1_f (new_AGEMA_signal_2086), .B0_t (key_s0_t[0]), .B0_f (key_s0_f[0]), .B1_t (key_s1_t[0]), .B1_f (key_s1_f[0]), .Z0_t (keyFF_MUX_inputPar_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_2090), .Z1_t (new_AGEMA_signal_2091), .Z1_f (new_AGEMA_signal_2092) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_2090), .B1_t (new_AGEMA_signal_2091), .B1_f (new_AGEMA_signal_2092), .Z0_t (keyFF_MUX_inputPar_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_2913), .Z1_t (new_AGEMA_signal_2914), .Z1_f (new_AGEMA_signal_2915) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_0_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_2913), .A1_t (new_AGEMA_signal_2914), .A1_f (new_AGEMA_signal_2915), .B0_t (keyFF_outputPar[3]), .B0_f (new_AGEMA_signal_2084), .B1_t (new_AGEMA_signal_2085), .B1_f (new_AGEMA_signal_2086), .Z0_t (keyFF_inputPar[0]), .Z0_f (new_AGEMA_signal_3373), .Z1_t (new_AGEMA_signal_3374), .Z1_f (new_AGEMA_signal_3375) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[4]), .A0_f (new_AGEMA_signal_2093), .A1_t (new_AGEMA_signal_2094), .A1_f (new_AGEMA_signal_2095), .B0_t (key_s0_t[1]), .B0_f (key_s0_f[1]), .B1_t (key_s1_t[1]), .B1_f (key_s1_f[1]), .Z0_t (keyFF_MUX_inputPar_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_2099), .Z1_t (new_AGEMA_signal_2100), .Z1_f (new_AGEMA_signal_2101) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_2099), .B1_t (new_AGEMA_signal_2100), .B1_f (new_AGEMA_signal_2101), .Z0_t (keyFF_MUX_inputPar_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_2916), .Z1_t (new_AGEMA_signal_2917), .Z1_f (new_AGEMA_signal_2918) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_1_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_2916), .A1_t (new_AGEMA_signal_2917), .A1_f (new_AGEMA_signal_2918), .B0_t (keyFF_outputPar[4]), .B0_f (new_AGEMA_signal_2093), .B1_t (new_AGEMA_signal_2094), .B1_f (new_AGEMA_signal_2095), .Z0_t (keyFF_inputPar[1]), .Z0_f (new_AGEMA_signal_3376), .Z1_t (new_AGEMA_signal_3377), .Z1_f (new_AGEMA_signal_3378) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[5]), .A0_f (new_AGEMA_signal_2102), .A1_t (new_AGEMA_signal_2103), .A1_f (new_AGEMA_signal_2104), .B0_t (key_s0_t[2]), .B0_f (key_s0_f[2]), .B1_t (key_s1_t[2]), .B1_f (key_s1_f[2]), .Z0_t (keyFF_MUX_inputPar_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_2108), .Z1_t (new_AGEMA_signal_2109), .Z1_f (new_AGEMA_signal_2110) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_2108), .B1_t (new_AGEMA_signal_2109), .B1_f (new_AGEMA_signal_2110), .Z0_t (keyFF_MUX_inputPar_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_2919), .Z1_t (new_AGEMA_signal_2920), .Z1_f (new_AGEMA_signal_2921) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_2_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_2919), .A1_t (new_AGEMA_signal_2920), .A1_f (new_AGEMA_signal_2921), .B0_t (keyFF_outputPar[5]), .B0_f (new_AGEMA_signal_2102), .B1_t (new_AGEMA_signal_2103), .B1_f (new_AGEMA_signal_2104), .Z0_t (keyFF_inputPar[2]), .Z0_f (new_AGEMA_signal_3379), .Z1_t (new_AGEMA_signal_3380), .Z1_f (new_AGEMA_signal_3381) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[6]), .A0_f (new_AGEMA_signal_2111), .A1_t (new_AGEMA_signal_2112), .A1_f (new_AGEMA_signal_2113), .B0_t (key_s0_t[3]), .B0_f (key_s0_f[3]), .B1_t (key_s1_t[3]), .B1_f (key_s1_f[3]), .Z0_t (keyFF_MUX_inputPar_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_2117), .Z1_t (new_AGEMA_signal_2118), .Z1_f (new_AGEMA_signal_2119) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_2117), .B1_t (new_AGEMA_signal_2118), .B1_f (new_AGEMA_signal_2119), .Z0_t (keyFF_MUX_inputPar_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_2922), .Z1_t (new_AGEMA_signal_2923), .Z1_f (new_AGEMA_signal_2924) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_3_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_2922), .A1_t (new_AGEMA_signal_2923), .A1_f (new_AGEMA_signal_2924), .B0_t (keyFF_outputPar[6]), .B0_f (new_AGEMA_signal_2111), .B1_t (new_AGEMA_signal_2112), .B1_f (new_AGEMA_signal_2113), .Z0_t (keyFF_inputPar[3]), .Z0_f (new_AGEMA_signal_3382), .Z1_t (new_AGEMA_signal_3383), .Z1_f (new_AGEMA_signal_3384) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[7]), .A0_f (new_AGEMA_signal_2120), .A1_t (new_AGEMA_signal_2121), .A1_f (new_AGEMA_signal_2122), .B0_t (key_s0_t[4]), .B0_f (key_s0_f[4]), .B1_t (key_s1_t[4]), .B1_f (key_s1_f[4]), .Z0_t (keyFF_MUX_inputPar_mux_inst_4_U1_X), .Z0_f (new_AGEMA_signal_2126), .Z1_t (new_AGEMA_signal_2127), .Z1_f (new_AGEMA_signal_2128) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_4_U1_X), .B0_f (new_AGEMA_signal_2126), .B1_t (new_AGEMA_signal_2127), .B1_f (new_AGEMA_signal_2128), .Z0_t (keyFF_MUX_inputPar_mux_inst_4_U1_Y), .Z0_f (new_AGEMA_signal_2925), .Z1_t (new_AGEMA_signal_2926), .Z1_f (new_AGEMA_signal_2927) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_4_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_4_U1_Y), .A0_f (new_AGEMA_signal_2925), .A1_t (new_AGEMA_signal_2926), .A1_f (new_AGEMA_signal_2927), .B0_t (keyFF_outputPar[7]), .B0_f (new_AGEMA_signal_2120), .B1_t (new_AGEMA_signal_2121), .B1_f (new_AGEMA_signal_2122), .Z0_t (keyFF_inputPar[4]), .Z0_f (new_AGEMA_signal_3385), .Z1_t (new_AGEMA_signal_3386), .Z1_f (new_AGEMA_signal_3387) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[8]), .A0_f (new_AGEMA_signal_2129), .A1_t (new_AGEMA_signal_2130), .A1_f (new_AGEMA_signal_2131), .B0_t (key_s0_t[5]), .B0_f (key_s0_f[5]), .B1_t (key_s1_t[5]), .B1_f (key_s1_f[5]), .Z0_t (keyFF_MUX_inputPar_mux_inst_5_U1_X), .Z0_f (new_AGEMA_signal_2135), .Z1_t (new_AGEMA_signal_2136), .Z1_f (new_AGEMA_signal_2137) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_5_U1_X), .B0_f (new_AGEMA_signal_2135), .B1_t (new_AGEMA_signal_2136), .B1_f (new_AGEMA_signal_2137), .Z0_t (keyFF_MUX_inputPar_mux_inst_5_U1_Y), .Z0_f (new_AGEMA_signal_2928), .Z1_t (new_AGEMA_signal_2929), .Z1_f (new_AGEMA_signal_2930) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_5_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_5_U1_Y), .A0_f (new_AGEMA_signal_2928), .A1_t (new_AGEMA_signal_2929), .A1_f (new_AGEMA_signal_2930), .B0_t (keyFF_outputPar[8]), .B0_f (new_AGEMA_signal_2129), .B1_t (new_AGEMA_signal_2130), .B1_f (new_AGEMA_signal_2131), .Z0_t (keyFF_inputPar[5]), .Z0_f (new_AGEMA_signal_3388), .Z1_t (new_AGEMA_signal_3389), .Z1_f (new_AGEMA_signal_3390) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[9]), .A0_f (new_AGEMA_signal_2138), .A1_t (new_AGEMA_signal_2139), .A1_f (new_AGEMA_signal_2140), .B0_t (key_s0_t[6]), .B0_f (key_s0_f[6]), .B1_t (key_s1_t[6]), .B1_f (key_s1_f[6]), .Z0_t (keyFF_MUX_inputPar_mux_inst_6_U1_X), .Z0_f (new_AGEMA_signal_2144), .Z1_t (new_AGEMA_signal_2145), .Z1_f (new_AGEMA_signal_2146) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_6_U1_X), .B0_f (new_AGEMA_signal_2144), .B1_t (new_AGEMA_signal_2145), .B1_f (new_AGEMA_signal_2146), .Z0_t (keyFF_MUX_inputPar_mux_inst_6_U1_Y), .Z0_f (new_AGEMA_signal_2931), .Z1_t (new_AGEMA_signal_2932), .Z1_f (new_AGEMA_signal_2933) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_6_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_6_U1_Y), .A0_f (new_AGEMA_signal_2931), .A1_t (new_AGEMA_signal_2932), .A1_f (new_AGEMA_signal_2933), .B0_t (keyFF_outputPar[9]), .B0_f (new_AGEMA_signal_2138), .B1_t (new_AGEMA_signal_2139), .B1_f (new_AGEMA_signal_2140), .Z0_t (keyFF_inputPar[6]), .Z0_f (new_AGEMA_signal_3391), .Z1_t (new_AGEMA_signal_3392), .Z1_f (new_AGEMA_signal_3393) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[10]), .A0_f (new_AGEMA_signal_2147), .A1_t (new_AGEMA_signal_2148), .A1_f (new_AGEMA_signal_2149), .B0_t (key_s0_t[7]), .B0_f (key_s0_f[7]), .B1_t (key_s1_t[7]), .B1_f (key_s1_f[7]), .Z0_t (keyFF_MUX_inputPar_mux_inst_7_U1_X), .Z0_f (new_AGEMA_signal_2153), .Z1_t (new_AGEMA_signal_2154), .Z1_f (new_AGEMA_signal_2155) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_7_U1_X), .B0_f (new_AGEMA_signal_2153), .B1_t (new_AGEMA_signal_2154), .B1_f (new_AGEMA_signal_2155), .Z0_t (keyFF_MUX_inputPar_mux_inst_7_U1_Y), .Z0_f (new_AGEMA_signal_2934), .Z1_t (new_AGEMA_signal_2935), .Z1_f (new_AGEMA_signal_2936) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_7_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_7_U1_Y), .A0_f (new_AGEMA_signal_2934), .A1_t (new_AGEMA_signal_2935), .A1_f (new_AGEMA_signal_2936), .B0_t (keyFF_outputPar[10]), .B0_f (new_AGEMA_signal_2147), .B1_t (new_AGEMA_signal_2148), .B1_f (new_AGEMA_signal_2149), .Z0_t (keyFF_inputPar[7]), .Z0_f (new_AGEMA_signal_3394), .Z1_t (new_AGEMA_signal_3395), .Z1_f (new_AGEMA_signal_3396) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[11]), .A0_f (new_AGEMA_signal_2156), .A1_t (new_AGEMA_signal_2157), .A1_f (new_AGEMA_signal_2158), .B0_t (key_s0_t[8]), .B0_f (key_s0_f[8]), .B1_t (key_s1_t[8]), .B1_f (key_s1_f[8]), .Z0_t (keyFF_MUX_inputPar_mux_inst_8_U1_X), .Z0_f (new_AGEMA_signal_2162), .Z1_t (new_AGEMA_signal_2163), .Z1_f (new_AGEMA_signal_2164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_8_U1_X), .B0_f (new_AGEMA_signal_2162), .B1_t (new_AGEMA_signal_2163), .B1_f (new_AGEMA_signal_2164), .Z0_t (keyFF_MUX_inputPar_mux_inst_8_U1_Y), .Z0_f (new_AGEMA_signal_2937), .Z1_t (new_AGEMA_signal_2938), .Z1_f (new_AGEMA_signal_2939) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_8_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_8_U1_Y), .A0_f (new_AGEMA_signal_2937), .A1_t (new_AGEMA_signal_2938), .A1_f (new_AGEMA_signal_2939), .B0_t (keyFF_outputPar[11]), .B0_f (new_AGEMA_signal_2156), .B1_t (new_AGEMA_signal_2157), .B1_f (new_AGEMA_signal_2158), .Z0_t (keyFF_inputPar[8]), .Z0_f (new_AGEMA_signal_3397), .Z1_t (new_AGEMA_signal_3398), .Z1_f (new_AGEMA_signal_3399) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[12]), .A0_f (new_AGEMA_signal_2165), .A1_t (new_AGEMA_signal_2166), .A1_f (new_AGEMA_signal_2167), .B0_t (key_s0_t[9]), .B0_f (key_s0_f[9]), .B1_t (key_s1_t[9]), .B1_f (key_s1_f[9]), .Z0_t (keyFF_MUX_inputPar_mux_inst_9_U1_X), .Z0_f (new_AGEMA_signal_2171), .Z1_t (new_AGEMA_signal_2172), .Z1_f (new_AGEMA_signal_2173) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_9_U1_X), .B0_f (new_AGEMA_signal_2171), .B1_t (new_AGEMA_signal_2172), .B1_f (new_AGEMA_signal_2173), .Z0_t (keyFF_MUX_inputPar_mux_inst_9_U1_Y), .Z0_f (new_AGEMA_signal_2940), .Z1_t (new_AGEMA_signal_2941), .Z1_f (new_AGEMA_signal_2942) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_9_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_9_U1_Y), .A0_f (new_AGEMA_signal_2940), .A1_t (new_AGEMA_signal_2941), .A1_f (new_AGEMA_signal_2942), .B0_t (keyFF_outputPar[12]), .B0_f (new_AGEMA_signal_2165), .B1_t (new_AGEMA_signal_2166), .B1_f (new_AGEMA_signal_2167), .Z0_t (keyFF_inputPar[9]), .Z0_f (new_AGEMA_signal_3400), .Z1_t (new_AGEMA_signal_3401), .Z1_f (new_AGEMA_signal_3402) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[13]), .A0_f (new_AGEMA_signal_2174), .A1_t (new_AGEMA_signal_2175), .A1_f (new_AGEMA_signal_2176), .B0_t (key_s0_t[10]), .B0_f (key_s0_f[10]), .B1_t (key_s1_t[10]), .B1_f (key_s1_f[10]), .Z0_t (keyFF_MUX_inputPar_mux_inst_10_U1_X), .Z0_f (new_AGEMA_signal_2180), .Z1_t (new_AGEMA_signal_2181), .Z1_f (new_AGEMA_signal_2182) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_10_U1_X), .B0_f (new_AGEMA_signal_2180), .B1_t (new_AGEMA_signal_2181), .B1_f (new_AGEMA_signal_2182), .Z0_t (keyFF_MUX_inputPar_mux_inst_10_U1_Y), .Z0_f (new_AGEMA_signal_2943), .Z1_t (new_AGEMA_signal_2944), .Z1_f (new_AGEMA_signal_2945) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_10_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_10_U1_Y), .A0_f (new_AGEMA_signal_2943), .A1_t (new_AGEMA_signal_2944), .A1_f (new_AGEMA_signal_2945), .B0_t (keyFF_outputPar[13]), .B0_f (new_AGEMA_signal_2174), .B1_t (new_AGEMA_signal_2175), .B1_f (new_AGEMA_signal_2176), .Z0_t (keyFF_inputPar[10]), .Z0_f (new_AGEMA_signal_3403), .Z1_t (new_AGEMA_signal_3404), .Z1_f (new_AGEMA_signal_3405) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[14]), .A0_f (new_AGEMA_signal_2183), .A1_t (new_AGEMA_signal_2184), .A1_f (new_AGEMA_signal_2185), .B0_t (key_s0_t[11]), .B0_f (key_s0_f[11]), .B1_t (key_s1_t[11]), .B1_f (key_s1_f[11]), .Z0_t (keyFF_MUX_inputPar_mux_inst_11_U1_X), .Z0_f (new_AGEMA_signal_2189), .Z1_t (new_AGEMA_signal_2190), .Z1_f (new_AGEMA_signal_2191) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_11_U1_X), .B0_f (new_AGEMA_signal_2189), .B1_t (new_AGEMA_signal_2190), .B1_f (new_AGEMA_signal_2191), .Z0_t (keyFF_MUX_inputPar_mux_inst_11_U1_Y), .Z0_f (new_AGEMA_signal_2946), .Z1_t (new_AGEMA_signal_2947), .Z1_f (new_AGEMA_signal_2948) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_11_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_11_U1_Y), .A0_f (new_AGEMA_signal_2946), .A1_t (new_AGEMA_signal_2947), .A1_f (new_AGEMA_signal_2948), .B0_t (keyFF_outputPar[14]), .B0_f (new_AGEMA_signal_2183), .B1_t (new_AGEMA_signal_2184), .B1_f (new_AGEMA_signal_2185), .Z0_t (keyFF_inputPar[11]), .Z0_f (new_AGEMA_signal_3406), .Z1_t (new_AGEMA_signal_3407), .Z1_f (new_AGEMA_signal_3408) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[15]), .A0_f (new_AGEMA_signal_2192), .A1_t (new_AGEMA_signal_2193), .A1_f (new_AGEMA_signal_2194), .B0_t (key_s0_t[12]), .B0_f (key_s0_f[12]), .B1_t (key_s1_t[12]), .B1_f (key_s1_f[12]), .Z0_t (keyFF_MUX_inputPar_mux_inst_12_U1_X), .Z0_f (new_AGEMA_signal_2198), .Z1_t (new_AGEMA_signal_2199), .Z1_f (new_AGEMA_signal_2200) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_12_U1_X), .B0_f (new_AGEMA_signal_2198), .B1_t (new_AGEMA_signal_2199), .B1_f (new_AGEMA_signal_2200), .Z0_t (keyFF_MUX_inputPar_mux_inst_12_U1_Y), .Z0_f (new_AGEMA_signal_2949), .Z1_t (new_AGEMA_signal_2950), .Z1_f (new_AGEMA_signal_2951) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_12_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_12_U1_Y), .A0_f (new_AGEMA_signal_2949), .A1_t (new_AGEMA_signal_2950), .A1_f (new_AGEMA_signal_2951), .B0_t (keyFF_outputPar[15]), .B0_f (new_AGEMA_signal_2192), .B1_t (new_AGEMA_signal_2193), .B1_f (new_AGEMA_signal_2194), .Z0_t (keyFF_inputPar[12]), .Z0_f (new_AGEMA_signal_3409), .Z1_t (new_AGEMA_signal_3410), .Z1_f (new_AGEMA_signal_3411) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[16]), .A0_f (new_AGEMA_signal_2201), .A1_t (new_AGEMA_signal_2202), .A1_f (new_AGEMA_signal_2203), .B0_t (key_s0_t[13]), .B0_f (key_s0_f[13]), .B1_t (key_s1_t[13]), .B1_f (key_s1_f[13]), .Z0_t (keyFF_MUX_inputPar_mux_inst_13_U1_X), .Z0_f (new_AGEMA_signal_2207), .Z1_t (new_AGEMA_signal_2208), .Z1_f (new_AGEMA_signal_2209) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_13_U1_X), .B0_f (new_AGEMA_signal_2207), .B1_t (new_AGEMA_signal_2208), .B1_f (new_AGEMA_signal_2209), .Z0_t (keyFF_MUX_inputPar_mux_inst_13_U1_Y), .Z0_f (new_AGEMA_signal_2952), .Z1_t (new_AGEMA_signal_2953), .Z1_f (new_AGEMA_signal_2954) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_13_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_13_U1_Y), .A0_f (new_AGEMA_signal_2952), .A1_t (new_AGEMA_signal_2953), .A1_f (new_AGEMA_signal_2954), .B0_t (keyFF_outputPar[16]), .B0_f (new_AGEMA_signal_2201), .B1_t (new_AGEMA_signal_2202), .B1_f (new_AGEMA_signal_2203), .Z0_t (keyFF_inputPar[13]), .Z0_f (new_AGEMA_signal_3412), .Z1_t (new_AGEMA_signal_3413), .Z1_f (new_AGEMA_signal_3414) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[17]), .A0_f (new_AGEMA_signal_2210), .A1_t (new_AGEMA_signal_2211), .A1_f (new_AGEMA_signal_2212), .B0_t (key_s0_t[14]), .B0_f (key_s0_f[14]), .B1_t (key_s1_t[14]), .B1_f (key_s1_f[14]), .Z0_t (keyFF_MUX_inputPar_mux_inst_14_U1_X), .Z0_f (new_AGEMA_signal_2216), .Z1_t (new_AGEMA_signal_2217), .Z1_f (new_AGEMA_signal_2218) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_14_U1_X), .B0_f (new_AGEMA_signal_2216), .B1_t (new_AGEMA_signal_2217), .B1_f (new_AGEMA_signal_2218), .Z0_t (keyFF_MUX_inputPar_mux_inst_14_U1_Y), .Z0_f (new_AGEMA_signal_2955), .Z1_t (new_AGEMA_signal_2956), .Z1_f (new_AGEMA_signal_2957) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_14_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_14_U1_Y), .A0_f (new_AGEMA_signal_2955), .A1_t (new_AGEMA_signal_2956), .A1_f (new_AGEMA_signal_2957), .B0_t (keyFF_outputPar[17]), .B0_f (new_AGEMA_signal_2210), .B1_t (new_AGEMA_signal_2211), .B1_f (new_AGEMA_signal_2212), .Z0_t (keyFF_inputPar[14]), .Z0_f (new_AGEMA_signal_3415), .Z1_t (new_AGEMA_signal_3416), .Z1_f (new_AGEMA_signal_3417) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[0]), .A0_f (new_AGEMA_signal_2075), .A1_t (new_AGEMA_signal_2076), .A1_f (new_AGEMA_signal_2077), .B0_t (key_s0_t[15]), .B0_f (key_s0_f[15]), .B1_t (key_s1_t[15]), .B1_f (key_s1_f[15]), .Z0_t (keyFF_MUX_inputPar_mux_inst_15_U1_X), .Z0_f (new_AGEMA_signal_2961), .Z1_t (new_AGEMA_signal_2962), .Z1_f (new_AGEMA_signal_2963) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_15_U1_X), .B0_f (new_AGEMA_signal_2961), .B1_t (new_AGEMA_signal_2962), .B1_f (new_AGEMA_signal_2963), .Z0_t (keyFF_MUX_inputPar_mux_inst_15_U1_Y), .Z0_f (new_AGEMA_signal_3418), .Z1_t (new_AGEMA_signal_3419), .Z1_f (new_AGEMA_signal_3420) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_15_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_15_U1_Y), .A0_f (new_AGEMA_signal_3418), .A1_t (new_AGEMA_signal_3419), .A1_f (new_AGEMA_signal_3420), .B0_t (keyFF_counterAdd[0]), .B0_f (new_AGEMA_signal_2075), .B1_t (new_AGEMA_signal_2076), .B1_f (new_AGEMA_signal_2077), .Z0_t (keyFF_inputPar[15]), .Z0_f (new_AGEMA_signal_4010), .Z1_t (new_AGEMA_signal_4011), .Z1_f (new_AGEMA_signal_4012) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[1]), .A0_f (new_AGEMA_signal_2063), .A1_t (new_AGEMA_signal_2064), .A1_f (new_AGEMA_signal_2065), .B0_t (key_s0_t[16]), .B0_f (key_s0_f[16]), .B1_t (key_s1_t[16]), .B1_f (key_s1_f[16]), .Z0_t (keyFF_MUX_inputPar_mux_inst_16_U1_X), .Z0_f (new_AGEMA_signal_2967), .Z1_t (new_AGEMA_signal_2968), .Z1_f (new_AGEMA_signal_2969) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_16_U1_X), .B0_f (new_AGEMA_signal_2967), .B1_t (new_AGEMA_signal_2968), .B1_f (new_AGEMA_signal_2969), .Z0_t (keyFF_MUX_inputPar_mux_inst_16_U1_Y), .Z0_f (new_AGEMA_signal_3421), .Z1_t (new_AGEMA_signal_3422), .Z1_f (new_AGEMA_signal_3423) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_16_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_16_U1_Y), .A0_f (new_AGEMA_signal_3421), .A1_t (new_AGEMA_signal_3422), .A1_f (new_AGEMA_signal_3423), .B0_t (keyFF_counterAdd[1]), .B0_f (new_AGEMA_signal_2063), .B1_t (new_AGEMA_signal_2064), .B1_f (new_AGEMA_signal_2065), .Z0_t (keyFF_inputPar[16]), .Z0_f (new_AGEMA_signal_4013), .Z1_t (new_AGEMA_signal_4014), .Z1_f (new_AGEMA_signal_4015) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[2]), .A0_f (new_AGEMA_signal_2081), .A1_t (new_AGEMA_signal_2082), .A1_f (new_AGEMA_signal_2083), .B0_t (key_s0_t[17]), .B0_f (key_s0_f[17]), .B1_t (key_s1_t[17]), .B1_f (key_s1_f[17]), .Z0_t (keyFF_MUX_inputPar_mux_inst_17_U1_X), .Z0_f (new_AGEMA_signal_2973), .Z1_t (new_AGEMA_signal_2974), .Z1_f (new_AGEMA_signal_2975) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_17_U1_X), .B0_f (new_AGEMA_signal_2973), .B1_t (new_AGEMA_signal_2974), .B1_f (new_AGEMA_signal_2975), .Z0_t (keyFF_MUX_inputPar_mux_inst_17_U1_Y), .Z0_f (new_AGEMA_signal_3424), .Z1_t (new_AGEMA_signal_3425), .Z1_f (new_AGEMA_signal_3426) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_17_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_17_U1_Y), .A0_f (new_AGEMA_signal_3424), .A1_t (new_AGEMA_signal_3425), .A1_f (new_AGEMA_signal_3426), .B0_t (keyFF_counterAdd[2]), .B0_f (new_AGEMA_signal_2081), .B1_t (new_AGEMA_signal_2082), .B1_f (new_AGEMA_signal_2083), .Z0_t (keyFF_inputPar[17]), .Z0_f (new_AGEMA_signal_4016), .Z1_t (new_AGEMA_signal_4017), .Z1_f (new_AGEMA_signal_4018) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[3]), .A0_f (new_AGEMA_signal_2057), .A1_t (new_AGEMA_signal_2058), .A1_f (new_AGEMA_signal_2059), .B0_t (key_s0_t[18]), .B0_f (key_s0_f[18]), .B1_t (key_s1_t[18]), .B1_f (key_s1_f[18]), .Z0_t (keyFF_MUX_inputPar_mux_inst_18_U1_X), .Z0_f (new_AGEMA_signal_2979), .Z1_t (new_AGEMA_signal_2980), .Z1_f (new_AGEMA_signal_2981) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_18_U1_X), .B0_f (new_AGEMA_signal_2979), .B1_t (new_AGEMA_signal_2980), .B1_f (new_AGEMA_signal_2981), .Z0_t (keyFF_MUX_inputPar_mux_inst_18_U1_Y), .Z0_f (new_AGEMA_signal_3427), .Z1_t (new_AGEMA_signal_3428), .Z1_f (new_AGEMA_signal_3429) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_18_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_18_U1_Y), .A0_f (new_AGEMA_signal_3427), .A1_t (new_AGEMA_signal_3428), .A1_f (new_AGEMA_signal_3429), .B0_t (keyFF_counterAdd[3]), .B0_f (new_AGEMA_signal_2057), .B1_t (new_AGEMA_signal_2058), .B1_f (new_AGEMA_signal_2059), .Z0_t (keyFF_inputPar[18]), .Z0_f (new_AGEMA_signal_4019), .Z1_t (new_AGEMA_signal_4020), .Z1_f (new_AGEMA_signal_4021) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_XOR1_U1 ( .A0_t (keyFF_counterAdd[4]), .A0_f (new_AGEMA_signal_2069), .A1_t (new_AGEMA_signal_2070), .A1_f (new_AGEMA_signal_2071), .B0_t (key_s0_t[19]), .B0_f (key_s0_f[19]), .B1_t (key_s1_t[19]), .B1_f (key_s1_f[19]), .Z0_t (keyFF_MUX_inputPar_mux_inst_19_U1_X), .Z0_f (new_AGEMA_signal_2985), .Z1_t (new_AGEMA_signal_2986), .Z1_f (new_AGEMA_signal_2987) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_19_U1_X), .B0_f (new_AGEMA_signal_2985), .B1_t (new_AGEMA_signal_2986), .B1_f (new_AGEMA_signal_2987), .Z0_t (keyFF_MUX_inputPar_mux_inst_19_U1_Y), .Z0_f (new_AGEMA_signal_3430), .Z1_t (new_AGEMA_signal_3431), .Z1_f (new_AGEMA_signal_3432) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_19_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_19_U1_Y), .A0_f (new_AGEMA_signal_3430), .A1_t (new_AGEMA_signal_3431), .A1_f (new_AGEMA_signal_3432), .B0_t (keyFF_counterAdd[4]), .B0_f (new_AGEMA_signal_2069), .B1_t (new_AGEMA_signal_2070), .B1_f (new_AGEMA_signal_2071), .Z0_t (keyFF_inputPar[19]), .Z0_f (new_AGEMA_signal_4022), .Z1_t (new_AGEMA_signal_4023), .Z1_f (new_AGEMA_signal_4024) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[23]), .A0_f (new_AGEMA_signal_2219), .A1_t (new_AGEMA_signal_2220), .A1_f (new_AGEMA_signal_2221), .B0_t (key_s0_t[20]), .B0_f (key_s0_f[20]), .B1_t (key_s1_t[20]), .B1_f (key_s1_f[20]), .Z0_t (keyFF_MUX_inputPar_mux_inst_20_U1_X), .Z0_f (new_AGEMA_signal_2225), .Z1_t (new_AGEMA_signal_2226), .Z1_f (new_AGEMA_signal_2227) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_20_U1_X), .B0_f (new_AGEMA_signal_2225), .B1_t (new_AGEMA_signal_2226), .B1_f (new_AGEMA_signal_2227), .Z0_t (keyFF_MUX_inputPar_mux_inst_20_U1_Y), .Z0_f (new_AGEMA_signal_2988), .Z1_t (new_AGEMA_signal_2989), .Z1_f (new_AGEMA_signal_2990) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_20_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_20_U1_Y), .A0_f (new_AGEMA_signal_2988), .A1_t (new_AGEMA_signal_2989), .A1_f (new_AGEMA_signal_2990), .B0_t (keyFF_outputPar[23]), .B0_f (new_AGEMA_signal_2219), .B1_t (new_AGEMA_signal_2220), .B1_f (new_AGEMA_signal_2221), .Z0_t (keyFF_inputPar[20]), .Z0_f (new_AGEMA_signal_3433), .Z1_t (new_AGEMA_signal_3434), .Z1_f (new_AGEMA_signal_3435) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[24]), .A0_f (new_AGEMA_signal_2228), .A1_t (new_AGEMA_signal_2229), .A1_f (new_AGEMA_signal_2230), .B0_t (key_s0_t[21]), .B0_f (key_s0_f[21]), .B1_t (key_s1_t[21]), .B1_f (key_s1_f[21]), .Z0_t (keyFF_MUX_inputPar_mux_inst_21_U1_X), .Z0_f (new_AGEMA_signal_2234), .Z1_t (new_AGEMA_signal_2235), .Z1_f (new_AGEMA_signal_2236) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_21_U1_X), .B0_f (new_AGEMA_signal_2234), .B1_t (new_AGEMA_signal_2235), .B1_f (new_AGEMA_signal_2236), .Z0_t (keyFF_MUX_inputPar_mux_inst_21_U1_Y), .Z0_f (new_AGEMA_signal_2991), .Z1_t (new_AGEMA_signal_2992), .Z1_f (new_AGEMA_signal_2993) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_21_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_21_U1_Y), .A0_f (new_AGEMA_signal_2991), .A1_t (new_AGEMA_signal_2992), .A1_f (new_AGEMA_signal_2993), .B0_t (keyFF_outputPar[24]), .B0_f (new_AGEMA_signal_2228), .B1_t (new_AGEMA_signal_2229), .B1_f (new_AGEMA_signal_2230), .Z0_t (keyFF_inputPar[21]), .Z0_f (new_AGEMA_signal_3436), .Z1_t (new_AGEMA_signal_3437), .Z1_f (new_AGEMA_signal_3438) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[25]), .A0_f (new_AGEMA_signal_2237), .A1_t (new_AGEMA_signal_2238), .A1_f (new_AGEMA_signal_2239), .B0_t (key_s0_t[22]), .B0_f (key_s0_f[22]), .B1_t (key_s1_t[22]), .B1_f (key_s1_f[22]), .Z0_t (keyFF_MUX_inputPar_mux_inst_22_U1_X), .Z0_f (new_AGEMA_signal_2243), .Z1_t (new_AGEMA_signal_2244), .Z1_f (new_AGEMA_signal_2245) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_22_U1_X), .B0_f (new_AGEMA_signal_2243), .B1_t (new_AGEMA_signal_2244), .B1_f (new_AGEMA_signal_2245), .Z0_t (keyFF_MUX_inputPar_mux_inst_22_U1_Y), .Z0_f (new_AGEMA_signal_2994), .Z1_t (new_AGEMA_signal_2995), .Z1_f (new_AGEMA_signal_2996) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_22_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_22_U1_Y), .A0_f (new_AGEMA_signal_2994), .A1_t (new_AGEMA_signal_2995), .A1_f (new_AGEMA_signal_2996), .B0_t (keyFF_outputPar[25]), .B0_f (new_AGEMA_signal_2237), .B1_t (new_AGEMA_signal_2238), .B1_f (new_AGEMA_signal_2239), .Z0_t (keyFF_inputPar[22]), .Z0_f (new_AGEMA_signal_3439), .Z1_t (new_AGEMA_signal_3440), .Z1_f (new_AGEMA_signal_3441) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[26]), .A0_f (new_AGEMA_signal_2246), .A1_t (new_AGEMA_signal_2247), .A1_f (new_AGEMA_signal_2248), .B0_t (key_s0_t[23]), .B0_f (key_s0_f[23]), .B1_t (key_s1_t[23]), .B1_f (key_s1_f[23]), .Z0_t (keyFF_MUX_inputPar_mux_inst_23_U1_X), .Z0_f (new_AGEMA_signal_2252), .Z1_t (new_AGEMA_signal_2253), .Z1_f (new_AGEMA_signal_2254) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_23_U1_X), .B0_f (new_AGEMA_signal_2252), .B1_t (new_AGEMA_signal_2253), .B1_f (new_AGEMA_signal_2254), .Z0_t (keyFF_MUX_inputPar_mux_inst_23_U1_Y), .Z0_f (new_AGEMA_signal_2997), .Z1_t (new_AGEMA_signal_2998), .Z1_f (new_AGEMA_signal_2999) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_23_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_23_U1_Y), .A0_f (new_AGEMA_signal_2997), .A1_t (new_AGEMA_signal_2998), .A1_f (new_AGEMA_signal_2999), .B0_t (keyFF_outputPar[26]), .B0_f (new_AGEMA_signal_2246), .B1_t (new_AGEMA_signal_2247), .B1_f (new_AGEMA_signal_2248), .Z0_t (keyFF_inputPar[23]), .Z0_f (new_AGEMA_signal_3442), .Z1_t (new_AGEMA_signal_3443), .Z1_f (new_AGEMA_signal_3444) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[27]), .A0_f (new_AGEMA_signal_2255), .A1_t (new_AGEMA_signal_2256), .A1_f (new_AGEMA_signal_2257), .B0_t (key_s0_t[24]), .B0_f (key_s0_f[24]), .B1_t (key_s1_t[24]), .B1_f (key_s1_f[24]), .Z0_t (keyFF_MUX_inputPar_mux_inst_24_U1_X), .Z0_f (new_AGEMA_signal_2261), .Z1_t (new_AGEMA_signal_2262), .Z1_f (new_AGEMA_signal_2263) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_24_U1_X), .B0_f (new_AGEMA_signal_2261), .B1_t (new_AGEMA_signal_2262), .B1_f (new_AGEMA_signal_2263), .Z0_t (keyFF_MUX_inputPar_mux_inst_24_U1_Y), .Z0_f (new_AGEMA_signal_3000), .Z1_t (new_AGEMA_signal_3001), .Z1_f (new_AGEMA_signal_3002) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_24_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_24_U1_Y), .A0_f (new_AGEMA_signal_3000), .A1_t (new_AGEMA_signal_3001), .A1_f (new_AGEMA_signal_3002), .B0_t (keyFF_outputPar[27]), .B0_f (new_AGEMA_signal_2255), .B1_t (new_AGEMA_signal_2256), .B1_f (new_AGEMA_signal_2257), .Z0_t (keyFF_inputPar[24]), .Z0_f (new_AGEMA_signal_3445), .Z1_t (new_AGEMA_signal_3446), .Z1_f (new_AGEMA_signal_3447) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[28]), .A0_f (new_AGEMA_signal_2264), .A1_t (new_AGEMA_signal_2265), .A1_f (new_AGEMA_signal_2266), .B0_t (key_s0_t[25]), .B0_f (key_s0_f[25]), .B1_t (key_s1_t[25]), .B1_f (key_s1_f[25]), .Z0_t (keyFF_MUX_inputPar_mux_inst_25_U1_X), .Z0_f (new_AGEMA_signal_2270), .Z1_t (new_AGEMA_signal_2271), .Z1_f (new_AGEMA_signal_2272) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_25_U1_X), .B0_f (new_AGEMA_signal_2270), .B1_t (new_AGEMA_signal_2271), .B1_f (new_AGEMA_signal_2272), .Z0_t (keyFF_MUX_inputPar_mux_inst_25_U1_Y), .Z0_f (new_AGEMA_signal_3003), .Z1_t (new_AGEMA_signal_3004), .Z1_f (new_AGEMA_signal_3005) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_25_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_25_U1_Y), .A0_f (new_AGEMA_signal_3003), .A1_t (new_AGEMA_signal_3004), .A1_f (new_AGEMA_signal_3005), .B0_t (keyFF_outputPar[28]), .B0_f (new_AGEMA_signal_2264), .B1_t (new_AGEMA_signal_2265), .B1_f (new_AGEMA_signal_2266), .Z0_t (keyFF_inputPar[25]), .Z0_f (new_AGEMA_signal_3448), .Z1_t (new_AGEMA_signal_3449), .Z1_f (new_AGEMA_signal_3450) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[29]), .A0_f (new_AGEMA_signal_2273), .A1_t (new_AGEMA_signal_2274), .A1_f (new_AGEMA_signal_2275), .B0_t (key_s0_t[26]), .B0_f (key_s0_f[26]), .B1_t (key_s1_t[26]), .B1_f (key_s1_f[26]), .Z0_t (keyFF_MUX_inputPar_mux_inst_26_U1_X), .Z0_f (new_AGEMA_signal_2279), .Z1_t (new_AGEMA_signal_2280), .Z1_f (new_AGEMA_signal_2281) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_26_U1_X), .B0_f (new_AGEMA_signal_2279), .B1_t (new_AGEMA_signal_2280), .B1_f (new_AGEMA_signal_2281), .Z0_t (keyFF_MUX_inputPar_mux_inst_26_U1_Y), .Z0_f (new_AGEMA_signal_3006), .Z1_t (new_AGEMA_signal_3007), .Z1_f (new_AGEMA_signal_3008) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_26_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_26_U1_Y), .A0_f (new_AGEMA_signal_3006), .A1_t (new_AGEMA_signal_3007), .A1_f (new_AGEMA_signal_3008), .B0_t (keyFF_outputPar[29]), .B0_f (new_AGEMA_signal_2273), .B1_t (new_AGEMA_signal_2274), .B1_f (new_AGEMA_signal_2275), .Z0_t (keyFF_inputPar[26]), .Z0_f (new_AGEMA_signal_3451), .Z1_t (new_AGEMA_signal_3452), .Z1_f (new_AGEMA_signal_3453) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[30]), .A0_f (new_AGEMA_signal_2282), .A1_t (new_AGEMA_signal_2283), .A1_f (new_AGEMA_signal_2284), .B0_t (key_s0_t[27]), .B0_f (key_s0_f[27]), .B1_t (key_s1_t[27]), .B1_f (key_s1_f[27]), .Z0_t (keyFF_MUX_inputPar_mux_inst_27_U1_X), .Z0_f (new_AGEMA_signal_2288), .Z1_t (new_AGEMA_signal_2289), .Z1_f (new_AGEMA_signal_2290) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_27_U1_X), .B0_f (new_AGEMA_signal_2288), .B1_t (new_AGEMA_signal_2289), .B1_f (new_AGEMA_signal_2290), .Z0_t (keyFF_MUX_inputPar_mux_inst_27_U1_Y), .Z0_f (new_AGEMA_signal_3009), .Z1_t (new_AGEMA_signal_3010), .Z1_f (new_AGEMA_signal_3011) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_27_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_27_U1_Y), .A0_f (new_AGEMA_signal_3009), .A1_t (new_AGEMA_signal_3010), .A1_f (new_AGEMA_signal_3011), .B0_t (keyFF_outputPar[30]), .B0_f (new_AGEMA_signal_2282), .B1_t (new_AGEMA_signal_2283), .B1_f (new_AGEMA_signal_2284), .Z0_t (keyFF_inputPar[27]), .Z0_f (new_AGEMA_signal_3454), .Z1_t (new_AGEMA_signal_3455), .Z1_f (new_AGEMA_signal_3456) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[31]), .A0_f (new_AGEMA_signal_2291), .A1_t (new_AGEMA_signal_2292), .A1_f (new_AGEMA_signal_2293), .B0_t (key_s0_t[28]), .B0_f (key_s0_f[28]), .B1_t (key_s1_t[28]), .B1_f (key_s1_f[28]), .Z0_t (keyFF_MUX_inputPar_mux_inst_28_U1_X), .Z0_f (new_AGEMA_signal_2297), .Z1_t (new_AGEMA_signal_2298), .Z1_f (new_AGEMA_signal_2299) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_28_U1_X), .B0_f (new_AGEMA_signal_2297), .B1_t (new_AGEMA_signal_2298), .B1_f (new_AGEMA_signal_2299), .Z0_t (keyFF_MUX_inputPar_mux_inst_28_U1_Y), .Z0_f (new_AGEMA_signal_3012), .Z1_t (new_AGEMA_signal_3013), .Z1_f (new_AGEMA_signal_3014) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_28_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_28_U1_Y), .A0_f (new_AGEMA_signal_3012), .A1_t (new_AGEMA_signal_3013), .A1_f (new_AGEMA_signal_3014), .B0_t (keyFF_outputPar[31]), .B0_f (new_AGEMA_signal_2291), .B1_t (new_AGEMA_signal_2292), .B1_f (new_AGEMA_signal_2293), .Z0_t (keyFF_inputPar[28]), .Z0_f (new_AGEMA_signal_3457), .Z1_t (new_AGEMA_signal_3458), .Z1_f (new_AGEMA_signal_3459) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[32]), .A0_f (new_AGEMA_signal_2300), .A1_t (new_AGEMA_signal_2301), .A1_f (new_AGEMA_signal_2302), .B0_t (key_s0_t[29]), .B0_f (key_s0_f[29]), .B1_t (key_s1_t[29]), .B1_f (key_s1_f[29]), .Z0_t (keyFF_MUX_inputPar_mux_inst_29_U1_X), .Z0_f (new_AGEMA_signal_2306), .Z1_t (new_AGEMA_signal_2307), .Z1_f (new_AGEMA_signal_2308) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_29_U1_X), .B0_f (new_AGEMA_signal_2306), .B1_t (new_AGEMA_signal_2307), .B1_f (new_AGEMA_signal_2308), .Z0_t (keyFF_MUX_inputPar_mux_inst_29_U1_Y), .Z0_f (new_AGEMA_signal_3015), .Z1_t (new_AGEMA_signal_3016), .Z1_f (new_AGEMA_signal_3017) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_29_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_29_U1_Y), .A0_f (new_AGEMA_signal_3015), .A1_t (new_AGEMA_signal_3016), .A1_f (new_AGEMA_signal_3017), .B0_t (keyFF_outputPar[32]), .B0_f (new_AGEMA_signal_2300), .B1_t (new_AGEMA_signal_2301), .B1_f (new_AGEMA_signal_2302), .Z0_t (keyFF_inputPar[29]), .Z0_f (new_AGEMA_signal_3460), .Z1_t (new_AGEMA_signal_3461), .Z1_f (new_AGEMA_signal_3462) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[33]), .A0_f (new_AGEMA_signal_2309), .A1_t (new_AGEMA_signal_2310), .A1_f (new_AGEMA_signal_2311), .B0_t (key_s0_t[30]), .B0_f (key_s0_f[30]), .B1_t (key_s1_t[30]), .B1_f (key_s1_f[30]), .Z0_t (keyFF_MUX_inputPar_mux_inst_30_U1_X), .Z0_f (new_AGEMA_signal_2315), .Z1_t (new_AGEMA_signal_2316), .Z1_f (new_AGEMA_signal_2317) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_30_U1_X), .B0_f (new_AGEMA_signal_2315), .B1_t (new_AGEMA_signal_2316), .B1_f (new_AGEMA_signal_2317), .Z0_t (keyFF_MUX_inputPar_mux_inst_30_U1_Y), .Z0_f (new_AGEMA_signal_3018), .Z1_t (new_AGEMA_signal_3019), .Z1_f (new_AGEMA_signal_3020) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_30_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_30_U1_Y), .A0_f (new_AGEMA_signal_3018), .A1_t (new_AGEMA_signal_3019), .A1_f (new_AGEMA_signal_3020), .B0_t (keyFF_outputPar[33]), .B0_f (new_AGEMA_signal_2309), .B1_t (new_AGEMA_signal_2310), .B1_f (new_AGEMA_signal_2311), .Z0_t (keyFF_inputPar[30]), .Z0_f (new_AGEMA_signal_3463), .Z1_t (new_AGEMA_signal_3464), .Z1_f (new_AGEMA_signal_3465) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[34]), .A0_f (new_AGEMA_signal_2318), .A1_t (new_AGEMA_signal_2319), .A1_f (new_AGEMA_signal_2320), .B0_t (key_s0_t[31]), .B0_f (key_s0_f[31]), .B1_t (key_s1_t[31]), .B1_f (key_s1_f[31]), .Z0_t (keyFF_MUX_inputPar_mux_inst_31_U1_X), .Z0_f (new_AGEMA_signal_2324), .Z1_t (new_AGEMA_signal_2325), .Z1_f (new_AGEMA_signal_2326) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_31_U1_X), .B0_f (new_AGEMA_signal_2324), .B1_t (new_AGEMA_signal_2325), .B1_f (new_AGEMA_signal_2326), .Z0_t (keyFF_MUX_inputPar_mux_inst_31_U1_Y), .Z0_f (new_AGEMA_signal_3021), .Z1_t (new_AGEMA_signal_3022), .Z1_f (new_AGEMA_signal_3023) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_31_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_31_U1_Y), .A0_f (new_AGEMA_signal_3021), .A1_t (new_AGEMA_signal_3022), .A1_f (new_AGEMA_signal_3023), .B0_t (keyFF_outputPar[34]), .B0_f (new_AGEMA_signal_2318), .B1_t (new_AGEMA_signal_2319), .B1_f (new_AGEMA_signal_2320), .Z0_t (keyFF_inputPar[31]), .Z0_f (new_AGEMA_signal_3466), .Z1_t (new_AGEMA_signal_3467), .Z1_f (new_AGEMA_signal_3468) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[35]), .A0_f (new_AGEMA_signal_2327), .A1_t (new_AGEMA_signal_2328), .A1_f (new_AGEMA_signal_2329), .B0_t (key_s0_t[32]), .B0_f (key_s0_f[32]), .B1_t (key_s1_t[32]), .B1_f (key_s1_f[32]), .Z0_t (keyFF_MUX_inputPar_mux_inst_32_U1_X), .Z0_f (new_AGEMA_signal_2333), .Z1_t (new_AGEMA_signal_2334), .Z1_f (new_AGEMA_signal_2335) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_32_U1_X), .B0_f (new_AGEMA_signal_2333), .B1_t (new_AGEMA_signal_2334), .B1_f (new_AGEMA_signal_2335), .Z0_t (keyFF_MUX_inputPar_mux_inst_32_U1_Y), .Z0_f (new_AGEMA_signal_3024), .Z1_t (new_AGEMA_signal_3025), .Z1_f (new_AGEMA_signal_3026) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_32_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_32_U1_Y), .A0_f (new_AGEMA_signal_3024), .A1_t (new_AGEMA_signal_3025), .A1_f (new_AGEMA_signal_3026), .B0_t (keyFF_outputPar[35]), .B0_f (new_AGEMA_signal_2327), .B1_t (new_AGEMA_signal_2328), .B1_f (new_AGEMA_signal_2329), .Z0_t (keyFF_inputPar[32]), .Z0_f (new_AGEMA_signal_3469), .Z1_t (new_AGEMA_signal_3470), .Z1_f (new_AGEMA_signal_3471) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[36]), .A0_f (new_AGEMA_signal_2336), .A1_t (new_AGEMA_signal_2337), .A1_f (new_AGEMA_signal_2338), .B0_t (key_s0_t[33]), .B0_f (key_s0_f[33]), .B1_t (key_s1_t[33]), .B1_f (key_s1_f[33]), .Z0_t (keyFF_MUX_inputPar_mux_inst_33_U1_X), .Z0_f (new_AGEMA_signal_2342), .Z1_t (new_AGEMA_signal_2343), .Z1_f (new_AGEMA_signal_2344) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_33_U1_X), .B0_f (new_AGEMA_signal_2342), .B1_t (new_AGEMA_signal_2343), .B1_f (new_AGEMA_signal_2344), .Z0_t (keyFF_MUX_inputPar_mux_inst_33_U1_Y), .Z0_f (new_AGEMA_signal_3027), .Z1_t (new_AGEMA_signal_3028), .Z1_f (new_AGEMA_signal_3029) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_33_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_33_U1_Y), .A0_f (new_AGEMA_signal_3027), .A1_t (new_AGEMA_signal_3028), .A1_f (new_AGEMA_signal_3029), .B0_t (keyFF_outputPar[36]), .B0_f (new_AGEMA_signal_2336), .B1_t (new_AGEMA_signal_2337), .B1_f (new_AGEMA_signal_2338), .Z0_t (keyFF_inputPar[33]), .Z0_f (new_AGEMA_signal_3472), .Z1_t (new_AGEMA_signal_3473), .Z1_f (new_AGEMA_signal_3474) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[37]), .A0_f (new_AGEMA_signal_2345), .A1_t (new_AGEMA_signal_2346), .A1_f (new_AGEMA_signal_2347), .B0_t (key_s0_t[34]), .B0_f (key_s0_f[34]), .B1_t (key_s1_t[34]), .B1_f (key_s1_f[34]), .Z0_t (keyFF_MUX_inputPar_mux_inst_34_U1_X), .Z0_f (new_AGEMA_signal_2351), .Z1_t (new_AGEMA_signal_2352), .Z1_f (new_AGEMA_signal_2353) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_34_U1_X), .B0_f (new_AGEMA_signal_2351), .B1_t (new_AGEMA_signal_2352), .B1_f (new_AGEMA_signal_2353), .Z0_t (keyFF_MUX_inputPar_mux_inst_34_U1_Y), .Z0_f (new_AGEMA_signal_3030), .Z1_t (new_AGEMA_signal_3031), .Z1_f (new_AGEMA_signal_3032) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_34_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_34_U1_Y), .A0_f (new_AGEMA_signal_3030), .A1_t (new_AGEMA_signal_3031), .A1_f (new_AGEMA_signal_3032), .B0_t (keyFF_outputPar[37]), .B0_f (new_AGEMA_signal_2345), .B1_t (new_AGEMA_signal_2346), .B1_f (new_AGEMA_signal_2347), .Z0_t (keyFF_inputPar[34]), .Z0_f (new_AGEMA_signal_3475), .Z1_t (new_AGEMA_signal_3476), .Z1_f (new_AGEMA_signal_3477) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[38]), .A0_f (new_AGEMA_signal_2354), .A1_t (new_AGEMA_signal_2355), .A1_f (new_AGEMA_signal_2356), .B0_t (key_s0_t[35]), .B0_f (key_s0_f[35]), .B1_t (key_s1_t[35]), .B1_f (key_s1_f[35]), .Z0_t (keyFF_MUX_inputPar_mux_inst_35_U1_X), .Z0_f (new_AGEMA_signal_2360), .Z1_t (new_AGEMA_signal_2361), .Z1_f (new_AGEMA_signal_2362) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_35_U1_X), .B0_f (new_AGEMA_signal_2360), .B1_t (new_AGEMA_signal_2361), .B1_f (new_AGEMA_signal_2362), .Z0_t (keyFF_MUX_inputPar_mux_inst_35_U1_Y), .Z0_f (new_AGEMA_signal_3033), .Z1_t (new_AGEMA_signal_3034), .Z1_f (new_AGEMA_signal_3035) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_35_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_35_U1_Y), .A0_f (new_AGEMA_signal_3033), .A1_t (new_AGEMA_signal_3034), .A1_f (new_AGEMA_signal_3035), .B0_t (keyFF_outputPar[38]), .B0_f (new_AGEMA_signal_2354), .B1_t (new_AGEMA_signal_2355), .B1_f (new_AGEMA_signal_2356), .Z0_t (keyFF_inputPar[35]), .Z0_f (new_AGEMA_signal_3478), .Z1_t (new_AGEMA_signal_3479), .Z1_f (new_AGEMA_signal_3480) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[39]), .A0_f (new_AGEMA_signal_2363), .A1_t (new_AGEMA_signal_2364), .A1_f (new_AGEMA_signal_2365), .B0_t (key_s0_t[36]), .B0_f (key_s0_f[36]), .B1_t (key_s1_t[36]), .B1_f (key_s1_f[36]), .Z0_t (keyFF_MUX_inputPar_mux_inst_36_U1_X), .Z0_f (new_AGEMA_signal_2369), .Z1_t (new_AGEMA_signal_2370), .Z1_f (new_AGEMA_signal_2371) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_36_U1_X), .B0_f (new_AGEMA_signal_2369), .B1_t (new_AGEMA_signal_2370), .B1_f (new_AGEMA_signal_2371), .Z0_t (keyFF_MUX_inputPar_mux_inst_36_U1_Y), .Z0_f (new_AGEMA_signal_3036), .Z1_t (new_AGEMA_signal_3037), .Z1_f (new_AGEMA_signal_3038) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_36_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_36_U1_Y), .A0_f (new_AGEMA_signal_3036), .A1_t (new_AGEMA_signal_3037), .A1_f (new_AGEMA_signal_3038), .B0_t (keyFF_outputPar[39]), .B0_f (new_AGEMA_signal_2363), .B1_t (new_AGEMA_signal_2364), .B1_f (new_AGEMA_signal_2365), .Z0_t (keyFF_inputPar[36]), .Z0_f (new_AGEMA_signal_3481), .Z1_t (new_AGEMA_signal_3482), .Z1_f (new_AGEMA_signal_3483) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[40]), .A0_f (new_AGEMA_signal_2372), .A1_t (new_AGEMA_signal_2373), .A1_f (new_AGEMA_signal_2374), .B0_t (key_s0_t[37]), .B0_f (key_s0_f[37]), .B1_t (key_s1_t[37]), .B1_f (key_s1_f[37]), .Z0_t (keyFF_MUX_inputPar_mux_inst_37_U1_X), .Z0_f (new_AGEMA_signal_2378), .Z1_t (new_AGEMA_signal_2379), .Z1_f (new_AGEMA_signal_2380) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_37_U1_X), .B0_f (new_AGEMA_signal_2378), .B1_t (new_AGEMA_signal_2379), .B1_f (new_AGEMA_signal_2380), .Z0_t (keyFF_MUX_inputPar_mux_inst_37_U1_Y), .Z0_f (new_AGEMA_signal_3039), .Z1_t (new_AGEMA_signal_3040), .Z1_f (new_AGEMA_signal_3041) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_37_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_37_U1_Y), .A0_f (new_AGEMA_signal_3039), .A1_t (new_AGEMA_signal_3040), .A1_f (new_AGEMA_signal_3041), .B0_t (keyFF_outputPar[40]), .B0_f (new_AGEMA_signal_2372), .B1_t (new_AGEMA_signal_2373), .B1_f (new_AGEMA_signal_2374), .Z0_t (keyFF_inputPar[37]), .Z0_f (new_AGEMA_signal_3484), .Z1_t (new_AGEMA_signal_3485), .Z1_f (new_AGEMA_signal_3486) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[41]), .A0_f (new_AGEMA_signal_2381), .A1_t (new_AGEMA_signal_2382), .A1_f (new_AGEMA_signal_2383), .B0_t (key_s0_t[38]), .B0_f (key_s0_f[38]), .B1_t (key_s1_t[38]), .B1_f (key_s1_f[38]), .Z0_t (keyFF_MUX_inputPar_mux_inst_38_U1_X), .Z0_f (new_AGEMA_signal_2387), .Z1_t (new_AGEMA_signal_2388), .Z1_f (new_AGEMA_signal_2389) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_38_U1_X), .B0_f (new_AGEMA_signal_2387), .B1_t (new_AGEMA_signal_2388), .B1_f (new_AGEMA_signal_2389), .Z0_t (keyFF_MUX_inputPar_mux_inst_38_U1_Y), .Z0_f (new_AGEMA_signal_3042), .Z1_t (new_AGEMA_signal_3043), .Z1_f (new_AGEMA_signal_3044) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_38_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_38_U1_Y), .A0_f (new_AGEMA_signal_3042), .A1_t (new_AGEMA_signal_3043), .A1_f (new_AGEMA_signal_3044), .B0_t (keyFF_outputPar[41]), .B0_f (new_AGEMA_signal_2381), .B1_t (new_AGEMA_signal_2382), .B1_f (new_AGEMA_signal_2383), .Z0_t (keyFF_inputPar[38]), .Z0_f (new_AGEMA_signal_3487), .Z1_t (new_AGEMA_signal_3488), .Z1_f (new_AGEMA_signal_3489) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[42]), .A0_f (new_AGEMA_signal_2390), .A1_t (new_AGEMA_signal_2391), .A1_f (new_AGEMA_signal_2392), .B0_t (key_s0_t[39]), .B0_f (key_s0_f[39]), .B1_t (key_s1_t[39]), .B1_f (key_s1_f[39]), .Z0_t (keyFF_MUX_inputPar_mux_inst_39_U1_X), .Z0_f (new_AGEMA_signal_2396), .Z1_t (new_AGEMA_signal_2397), .Z1_f (new_AGEMA_signal_2398) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_39_U1_X), .B0_f (new_AGEMA_signal_2396), .B1_t (new_AGEMA_signal_2397), .B1_f (new_AGEMA_signal_2398), .Z0_t (keyFF_MUX_inputPar_mux_inst_39_U1_Y), .Z0_f (new_AGEMA_signal_3045), .Z1_t (new_AGEMA_signal_3046), .Z1_f (new_AGEMA_signal_3047) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_39_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_39_U1_Y), .A0_f (new_AGEMA_signal_3045), .A1_t (new_AGEMA_signal_3046), .A1_f (new_AGEMA_signal_3047), .B0_t (keyFF_outputPar[42]), .B0_f (new_AGEMA_signal_2390), .B1_t (new_AGEMA_signal_2391), .B1_f (new_AGEMA_signal_2392), .Z0_t (keyFF_inputPar[39]), .Z0_f (new_AGEMA_signal_3490), .Z1_t (new_AGEMA_signal_3491), .Z1_f (new_AGEMA_signal_3492) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[43]), .A0_f (new_AGEMA_signal_2399), .A1_t (new_AGEMA_signal_2400), .A1_f (new_AGEMA_signal_2401), .B0_t (key_s0_t[40]), .B0_f (key_s0_f[40]), .B1_t (key_s1_t[40]), .B1_f (key_s1_f[40]), .Z0_t (keyFF_MUX_inputPar_mux_inst_40_U1_X), .Z0_f (new_AGEMA_signal_2405), .Z1_t (new_AGEMA_signal_2406), .Z1_f (new_AGEMA_signal_2407) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_40_U1_X), .B0_f (new_AGEMA_signal_2405), .B1_t (new_AGEMA_signal_2406), .B1_f (new_AGEMA_signal_2407), .Z0_t (keyFF_MUX_inputPar_mux_inst_40_U1_Y), .Z0_f (new_AGEMA_signal_3048), .Z1_t (new_AGEMA_signal_3049), .Z1_f (new_AGEMA_signal_3050) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_40_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_40_U1_Y), .A0_f (new_AGEMA_signal_3048), .A1_t (new_AGEMA_signal_3049), .A1_f (new_AGEMA_signal_3050), .B0_t (keyFF_outputPar[43]), .B0_f (new_AGEMA_signal_2399), .B1_t (new_AGEMA_signal_2400), .B1_f (new_AGEMA_signal_2401), .Z0_t (keyFF_inputPar[40]), .Z0_f (new_AGEMA_signal_3493), .Z1_t (new_AGEMA_signal_3494), .Z1_f (new_AGEMA_signal_3495) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[44]), .A0_f (new_AGEMA_signal_2408), .A1_t (new_AGEMA_signal_2409), .A1_f (new_AGEMA_signal_2410), .B0_t (key_s0_t[41]), .B0_f (key_s0_f[41]), .B1_t (key_s1_t[41]), .B1_f (key_s1_f[41]), .Z0_t (keyFF_MUX_inputPar_mux_inst_41_U1_X), .Z0_f (new_AGEMA_signal_2414), .Z1_t (new_AGEMA_signal_2415), .Z1_f (new_AGEMA_signal_2416) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_41_U1_X), .B0_f (new_AGEMA_signal_2414), .B1_t (new_AGEMA_signal_2415), .B1_f (new_AGEMA_signal_2416), .Z0_t (keyFF_MUX_inputPar_mux_inst_41_U1_Y), .Z0_f (new_AGEMA_signal_3051), .Z1_t (new_AGEMA_signal_3052), .Z1_f (new_AGEMA_signal_3053) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_41_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_41_U1_Y), .A0_f (new_AGEMA_signal_3051), .A1_t (new_AGEMA_signal_3052), .A1_f (new_AGEMA_signal_3053), .B0_t (keyFF_outputPar[44]), .B0_f (new_AGEMA_signal_2408), .B1_t (new_AGEMA_signal_2409), .B1_f (new_AGEMA_signal_2410), .Z0_t (keyFF_inputPar[41]), .Z0_f (new_AGEMA_signal_3496), .Z1_t (new_AGEMA_signal_3497), .Z1_f (new_AGEMA_signal_3498) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[45]), .A0_f (new_AGEMA_signal_2417), .A1_t (new_AGEMA_signal_2418), .A1_f (new_AGEMA_signal_2419), .B0_t (key_s0_t[42]), .B0_f (key_s0_f[42]), .B1_t (key_s1_t[42]), .B1_f (key_s1_f[42]), .Z0_t (keyFF_MUX_inputPar_mux_inst_42_U1_X), .Z0_f (new_AGEMA_signal_2423), .Z1_t (new_AGEMA_signal_2424), .Z1_f (new_AGEMA_signal_2425) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_42_U1_X), .B0_f (new_AGEMA_signal_2423), .B1_t (new_AGEMA_signal_2424), .B1_f (new_AGEMA_signal_2425), .Z0_t (keyFF_MUX_inputPar_mux_inst_42_U1_Y), .Z0_f (new_AGEMA_signal_3054), .Z1_t (new_AGEMA_signal_3055), .Z1_f (new_AGEMA_signal_3056) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_42_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_42_U1_Y), .A0_f (new_AGEMA_signal_3054), .A1_t (new_AGEMA_signal_3055), .A1_f (new_AGEMA_signal_3056), .B0_t (keyFF_outputPar[45]), .B0_f (new_AGEMA_signal_2417), .B1_t (new_AGEMA_signal_2418), .B1_f (new_AGEMA_signal_2419), .Z0_t (keyFF_inputPar[42]), .Z0_f (new_AGEMA_signal_3499), .Z1_t (new_AGEMA_signal_3500), .Z1_f (new_AGEMA_signal_3501) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[46]), .A0_f (new_AGEMA_signal_2426), .A1_t (new_AGEMA_signal_2427), .A1_f (new_AGEMA_signal_2428), .B0_t (key_s0_t[43]), .B0_f (key_s0_f[43]), .B1_t (key_s1_t[43]), .B1_f (key_s1_f[43]), .Z0_t (keyFF_MUX_inputPar_mux_inst_43_U1_X), .Z0_f (new_AGEMA_signal_2432), .Z1_t (new_AGEMA_signal_2433), .Z1_f (new_AGEMA_signal_2434) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_43_U1_X), .B0_f (new_AGEMA_signal_2432), .B1_t (new_AGEMA_signal_2433), .B1_f (new_AGEMA_signal_2434), .Z0_t (keyFF_MUX_inputPar_mux_inst_43_U1_Y), .Z0_f (new_AGEMA_signal_3057), .Z1_t (new_AGEMA_signal_3058), .Z1_f (new_AGEMA_signal_3059) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_43_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_43_U1_Y), .A0_f (new_AGEMA_signal_3057), .A1_t (new_AGEMA_signal_3058), .A1_f (new_AGEMA_signal_3059), .B0_t (keyFF_outputPar[46]), .B0_f (new_AGEMA_signal_2426), .B1_t (new_AGEMA_signal_2427), .B1_f (new_AGEMA_signal_2428), .Z0_t (keyFF_inputPar[43]), .Z0_f (new_AGEMA_signal_3502), .Z1_t (new_AGEMA_signal_3503), .Z1_f (new_AGEMA_signal_3504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[47]), .A0_f (new_AGEMA_signal_2435), .A1_t (new_AGEMA_signal_2436), .A1_f (new_AGEMA_signal_2437), .B0_t (key_s0_t[44]), .B0_f (key_s0_f[44]), .B1_t (key_s1_t[44]), .B1_f (key_s1_f[44]), .Z0_t (keyFF_MUX_inputPar_mux_inst_44_U1_X), .Z0_f (new_AGEMA_signal_2441), .Z1_t (new_AGEMA_signal_2442), .Z1_f (new_AGEMA_signal_2443) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_44_U1_X), .B0_f (new_AGEMA_signal_2441), .B1_t (new_AGEMA_signal_2442), .B1_f (new_AGEMA_signal_2443), .Z0_t (keyFF_MUX_inputPar_mux_inst_44_U1_Y), .Z0_f (new_AGEMA_signal_3060), .Z1_t (new_AGEMA_signal_3061), .Z1_f (new_AGEMA_signal_3062) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_44_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_44_U1_Y), .A0_f (new_AGEMA_signal_3060), .A1_t (new_AGEMA_signal_3061), .A1_f (new_AGEMA_signal_3062), .B0_t (keyFF_outputPar[47]), .B0_f (new_AGEMA_signal_2435), .B1_t (new_AGEMA_signal_2436), .B1_f (new_AGEMA_signal_2437), .Z0_t (keyFF_inputPar[44]), .Z0_f (new_AGEMA_signal_3505), .Z1_t (new_AGEMA_signal_3506), .Z1_f (new_AGEMA_signal_3507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[48]), .A0_f (new_AGEMA_signal_2444), .A1_t (new_AGEMA_signal_2445), .A1_f (new_AGEMA_signal_2446), .B0_t (key_s0_t[45]), .B0_f (key_s0_f[45]), .B1_t (key_s1_t[45]), .B1_f (key_s1_f[45]), .Z0_t (keyFF_MUX_inputPar_mux_inst_45_U1_X), .Z0_f (new_AGEMA_signal_2450), .Z1_t (new_AGEMA_signal_2451), .Z1_f (new_AGEMA_signal_2452) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_45_U1_X), .B0_f (new_AGEMA_signal_2450), .B1_t (new_AGEMA_signal_2451), .B1_f (new_AGEMA_signal_2452), .Z0_t (keyFF_MUX_inputPar_mux_inst_45_U1_Y), .Z0_f (new_AGEMA_signal_3063), .Z1_t (new_AGEMA_signal_3064), .Z1_f (new_AGEMA_signal_3065) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_45_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_45_U1_Y), .A0_f (new_AGEMA_signal_3063), .A1_t (new_AGEMA_signal_3064), .A1_f (new_AGEMA_signal_3065), .B0_t (keyFF_outputPar[48]), .B0_f (new_AGEMA_signal_2444), .B1_t (new_AGEMA_signal_2445), .B1_f (new_AGEMA_signal_2446), .Z0_t (keyFF_inputPar[45]), .Z0_f (new_AGEMA_signal_3508), .Z1_t (new_AGEMA_signal_3509), .Z1_f (new_AGEMA_signal_3510) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[49]), .A0_f (new_AGEMA_signal_2453), .A1_t (new_AGEMA_signal_2454), .A1_f (new_AGEMA_signal_2455), .B0_t (key_s0_t[46]), .B0_f (key_s0_f[46]), .B1_t (key_s1_t[46]), .B1_f (key_s1_f[46]), .Z0_t (keyFF_MUX_inputPar_mux_inst_46_U1_X), .Z0_f (new_AGEMA_signal_2459), .Z1_t (new_AGEMA_signal_2460), .Z1_f (new_AGEMA_signal_2461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_46_U1_X), .B0_f (new_AGEMA_signal_2459), .B1_t (new_AGEMA_signal_2460), .B1_f (new_AGEMA_signal_2461), .Z0_t (keyFF_MUX_inputPar_mux_inst_46_U1_Y), .Z0_f (new_AGEMA_signal_3066), .Z1_t (new_AGEMA_signal_3067), .Z1_f (new_AGEMA_signal_3068) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_46_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_46_U1_Y), .A0_f (new_AGEMA_signal_3066), .A1_t (new_AGEMA_signal_3067), .A1_f (new_AGEMA_signal_3068), .B0_t (keyFF_outputPar[49]), .B0_f (new_AGEMA_signal_2453), .B1_t (new_AGEMA_signal_2454), .B1_f (new_AGEMA_signal_2455), .Z0_t (keyFF_inputPar[46]), .Z0_f (new_AGEMA_signal_3511), .Z1_t (new_AGEMA_signal_3512), .Z1_f (new_AGEMA_signal_3513) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[50]), .A0_f (new_AGEMA_signal_2462), .A1_t (new_AGEMA_signal_2463), .A1_f (new_AGEMA_signal_2464), .B0_t (key_s0_t[47]), .B0_f (key_s0_f[47]), .B1_t (key_s1_t[47]), .B1_f (key_s1_f[47]), .Z0_t (keyFF_MUX_inputPar_mux_inst_47_U1_X), .Z0_f (new_AGEMA_signal_2468), .Z1_t (new_AGEMA_signal_2469), .Z1_f (new_AGEMA_signal_2470) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_47_U1_X), .B0_f (new_AGEMA_signal_2468), .B1_t (new_AGEMA_signal_2469), .B1_f (new_AGEMA_signal_2470), .Z0_t (keyFF_MUX_inputPar_mux_inst_47_U1_Y), .Z0_f (new_AGEMA_signal_3069), .Z1_t (new_AGEMA_signal_3070), .Z1_f (new_AGEMA_signal_3071) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_47_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_47_U1_Y), .A0_f (new_AGEMA_signal_3069), .A1_t (new_AGEMA_signal_3070), .A1_f (new_AGEMA_signal_3071), .B0_t (keyFF_outputPar[50]), .B0_f (new_AGEMA_signal_2462), .B1_t (new_AGEMA_signal_2463), .B1_f (new_AGEMA_signal_2464), .Z0_t (keyFF_inputPar[47]), .Z0_f (new_AGEMA_signal_3514), .Z1_t (new_AGEMA_signal_3515), .Z1_f (new_AGEMA_signal_3516) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[51]), .A0_f (new_AGEMA_signal_2471), .A1_t (new_AGEMA_signal_2472), .A1_f (new_AGEMA_signal_2473), .B0_t (key_s0_t[48]), .B0_f (key_s0_f[48]), .B1_t (key_s1_t[48]), .B1_f (key_s1_f[48]), .Z0_t (keyFF_MUX_inputPar_mux_inst_48_U1_X), .Z0_f (new_AGEMA_signal_2477), .Z1_t (new_AGEMA_signal_2478), .Z1_f (new_AGEMA_signal_2479) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_48_U1_X), .B0_f (new_AGEMA_signal_2477), .B1_t (new_AGEMA_signal_2478), .B1_f (new_AGEMA_signal_2479), .Z0_t (keyFF_MUX_inputPar_mux_inst_48_U1_Y), .Z0_f (new_AGEMA_signal_3072), .Z1_t (new_AGEMA_signal_3073), .Z1_f (new_AGEMA_signal_3074) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_48_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_48_U1_Y), .A0_f (new_AGEMA_signal_3072), .A1_t (new_AGEMA_signal_3073), .A1_f (new_AGEMA_signal_3074), .B0_t (keyFF_outputPar[51]), .B0_f (new_AGEMA_signal_2471), .B1_t (new_AGEMA_signal_2472), .B1_f (new_AGEMA_signal_2473), .Z0_t (keyFF_inputPar[48]), .Z0_f (new_AGEMA_signal_3517), .Z1_t (new_AGEMA_signal_3518), .Z1_f (new_AGEMA_signal_3519) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[52]), .A0_f (new_AGEMA_signal_2480), .A1_t (new_AGEMA_signal_2481), .A1_f (new_AGEMA_signal_2482), .B0_t (key_s0_t[49]), .B0_f (key_s0_f[49]), .B1_t (key_s1_t[49]), .B1_f (key_s1_f[49]), .Z0_t (keyFF_MUX_inputPar_mux_inst_49_U1_X), .Z0_f (new_AGEMA_signal_2486), .Z1_t (new_AGEMA_signal_2487), .Z1_f (new_AGEMA_signal_2488) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_49_U1_X), .B0_f (new_AGEMA_signal_2486), .B1_t (new_AGEMA_signal_2487), .B1_f (new_AGEMA_signal_2488), .Z0_t (keyFF_MUX_inputPar_mux_inst_49_U1_Y), .Z0_f (new_AGEMA_signal_3075), .Z1_t (new_AGEMA_signal_3076), .Z1_f (new_AGEMA_signal_3077) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_49_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_49_U1_Y), .A0_f (new_AGEMA_signal_3075), .A1_t (new_AGEMA_signal_3076), .A1_f (new_AGEMA_signal_3077), .B0_t (keyFF_outputPar[52]), .B0_f (new_AGEMA_signal_2480), .B1_t (new_AGEMA_signal_2481), .B1_f (new_AGEMA_signal_2482), .Z0_t (keyFF_inputPar[49]), .Z0_f (new_AGEMA_signal_3520), .Z1_t (new_AGEMA_signal_3521), .Z1_f (new_AGEMA_signal_3522) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[53]), .A0_f (new_AGEMA_signal_2489), .A1_t (new_AGEMA_signal_2490), .A1_f (new_AGEMA_signal_2491), .B0_t (key_s0_t[50]), .B0_f (key_s0_f[50]), .B1_t (key_s1_t[50]), .B1_f (key_s1_f[50]), .Z0_t (keyFF_MUX_inputPar_mux_inst_50_U1_X), .Z0_f (new_AGEMA_signal_2495), .Z1_t (new_AGEMA_signal_2496), .Z1_f (new_AGEMA_signal_2497) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_50_U1_X), .B0_f (new_AGEMA_signal_2495), .B1_t (new_AGEMA_signal_2496), .B1_f (new_AGEMA_signal_2497), .Z0_t (keyFF_MUX_inputPar_mux_inst_50_U1_Y), .Z0_f (new_AGEMA_signal_3078), .Z1_t (new_AGEMA_signal_3079), .Z1_f (new_AGEMA_signal_3080) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_50_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_50_U1_Y), .A0_f (new_AGEMA_signal_3078), .A1_t (new_AGEMA_signal_3079), .A1_f (new_AGEMA_signal_3080), .B0_t (keyFF_outputPar[53]), .B0_f (new_AGEMA_signal_2489), .B1_t (new_AGEMA_signal_2490), .B1_f (new_AGEMA_signal_2491), .Z0_t (keyFF_inputPar[50]), .Z0_f (new_AGEMA_signal_3523), .Z1_t (new_AGEMA_signal_3524), .Z1_f (new_AGEMA_signal_3525) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[54]), .A0_f (new_AGEMA_signal_2498), .A1_t (new_AGEMA_signal_2499), .A1_f (new_AGEMA_signal_2500), .B0_t (key_s0_t[51]), .B0_f (key_s0_f[51]), .B1_t (key_s1_t[51]), .B1_f (key_s1_f[51]), .Z0_t (keyFF_MUX_inputPar_mux_inst_51_U1_X), .Z0_f (new_AGEMA_signal_2504), .Z1_t (new_AGEMA_signal_2505), .Z1_f (new_AGEMA_signal_2506) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_51_U1_X), .B0_f (new_AGEMA_signal_2504), .B1_t (new_AGEMA_signal_2505), .B1_f (new_AGEMA_signal_2506), .Z0_t (keyFF_MUX_inputPar_mux_inst_51_U1_Y), .Z0_f (new_AGEMA_signal_3081), .Z1_t (new_AGEMA_signal_3082), .Z1_f (new_AGEMA_signal_3083) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_51_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_51_U1_Y), .A0_f (new_AGEMA_signal_3081), .A1_t (new_AGEMA_signal_3082), .A1_f (new_AGEMA_signal_3083), .B0_t (keyFF_outputPar[54]), .B0_f (new_AGEMA_signal_2498), .B1_t (new_AGEMA_signal_2499), .B1_f (new_AGEMA_signal_2500), .Z0_t (keyFF_inputPar[51]), .Z0_f (new_AGEMA_signal_3526), .Z1_t (new_AGEMA_signal_3527), .Z1_f (new_AGEMA_signal_3528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[55]), .A0_f (new_AGEMA_signal_2507), .A1_t (new_AGEMA_signal_2508), .A1_f (new_AGEMA_signal_2509), .B0_t (key_s0_t[52]), .B0_f (key_s0_f[52]), .B1_t (key_s1_t[52]), .B1_f (key_s1_f[52]), .Z0_t (keyFF_MUX_inputPar_mux_inst_52_U1_X), .Z0_f (new_AGEMA_signal_2513), .Z1_t (new_AGEMA_signal_2514), .Z1_f (new_AGEMA_signal_2515) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_52_U1_X), .B0_f (new_AGEMA_signal_2513), .B1_t (new_AGEMA_signal_2514), .B1_f (new_AGEMA_signal_2515), .Z0_t (keyFF_MUX_inputPar_mux_inst_52_U1_Y), .Z0_f (new_AGEMA_signal_3084), .Z1_t (new_AGEMA_signal_3085), .Z1_f (new_AGEMA_signal_3086) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_52_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_52_U1_Y), .A0_f (new_AGEMA_signal_3084), .A1_t (new_AGEMA_signal_3085), .A1_f (new_AGEMA_signal_3086), .B0_t (keyFF_outputPar[55]), .B0_f (new_AGEMA_signal_2507), .B1_t (new_AGEMA_signal_2508), .B1_f (new_AGEMA_signal_2509), .Z0_t (keyFF_inputPar[52]), .Z0_f (new_AGEMA_signal_3529), .Z1_t (new_AGEMA_signal_3530), .Z1_f (new_AGEMA_signal_3531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[56]), .A0_f (new_AGEMA_signal_2516), .A1_t (new_AGEMA_signal_2517), .A1_f (new_AGEMA_signal_2518), .B0_t (key_s0_t[53]), .B0_f (key_s0_f[53]), .B1_t (key_s1_t[53]), .B1_f (key_s1_f[53]), .Z0_t (keyFF_MUX_inputPar_mux_inst_53_U1_X), .Z0_f (new_AGEMA_signal_2522), .Z1_t (new_AGEMA_signal_2523), .Z1_f (new_AGEMA_signal_2524) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_53_U1_X), .B0_f (new_AGEMA_signal_2522), .B1_t (new_AGEMA_signal_2523), .B1_f (new_AGEMA_signal_2524), .Z0_t (keyFF_MUX_inputPar_mux_inst_53_U1_Y), .Z0_f (new_AGEMA_signal_3087), .Z1_t (new_AGEMA_signal_3088), .Z1_f (new_AGEMA_signal_3089) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_53_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_53_U1_Y), .A0_f (new_AGEMA_signal_3087), .A1_t (new_AGEMA_signal_3088), .A1_f (new_AGEMA_signal_3089), .B0_t (keyFF_outputPar[56]), .B0_f (new_AGEMA_signal_2516), .B1_t (new_AGEMA_signal_2517), .B1_f (new_AGEMA_signal_2518), .Z0_t (keyFF_inputPar[53]), .Z0_f (new_AGEMA_signal_3532), .Z1_t (new_AGEMA_signal_3533), .Z1_f (new_AGEMA_signal_3534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[57]), .A0_f (new_AGEMA_signal_2525), .A1_t (new_AGEMA_signal_2526), .A1_f (new_AGEMA_signal_2527), .B0_t (key_s0_t[54]), .B0_f (key_s0_f[54]), .B1_t (key_s1_t[54]), .B1_f (key_s1_f[54]), .Z0_t (keyFF_MUX_inputPar_mux_inst_54_U1_X), .Z0_f (new_AGEMA_signal_2531), .Z1_t (new_AGEMA_signal_2532), .Z1_f (new_AGEMA_signal_2533) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_54_U1_X), .B0_f (new_AGEMA_signal_2531), .B1_t (new_AGEMA_signal_2532), .B1_f (new_AGEMA_signal_2533), .Z0_t (keyFF_MUX_inputPar_mux_inst_54_U1_Y), .Z0_f (new_AGEMA_signal_3090), .Z1_t (new_AGEMA_signal_3091), .Z1_f (new_AGEMA_signal_3092) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_54_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_54_U1_Y), .A0_f (new_AGEMA_signal_3090), .A1_t (new_AGEMA_signal_3091), .A1_f (new_AGEMA_signal_3092), .B0_t (keyFF_outputPar[57]), .B0_f (new_AGEMA_signal_2525), .B1_t (new_AGEMA_signal_2526), .B1_f (new_AGEMA_signal_2527), .Z0_t (keyFF_inputPar[54]), .Z0_f (new_AGEMA_signal_3535), .Z1_t (new_AGEMA_signal_3536), .Z1_f (new_AGEMA_signal_3537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[58]), .A0_f (new_AGEMA_signal_2534), .A1_t (new_AGEMA_signal_2535), .A1_f (new_AGEMA_signal_2536), .B0_t (key_s0_t[55]), .B0_f (key_s0_f[55]), .B1_t (key_s1_t[55]), .B1_f (key_s1_f[55]), .Z0_t (keyFF_MUX_inputPar_mux_inst_55_U1_X), .Z0_f (new_AGEMA_signal_2540), .Z1_t (new_AGEMA_signal_2541), .Z1_f (new_AGEMA_signal_2542) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_55_U1_X), .B0_f (new_AGEMA_signal_2540), .B1_t (new_AGEMA_signal_2541), .B1_f (new_AGEMA_signal_2542), .Z0_t (keyFF_MUX_inputPar_mux_inst_55_U1_Y), .Z0_f (new_AGEMA_signal_3093), .Z1_t (new_AGEMA_signal_3094), .Z1_f (new_AGEMA_signal_3095) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_55_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_55_U1_Y), .A0_f (new_AGEMA_signal_3093), .A1_t (new_AGEMA_signal_3094), .A1_f (new_AGEMA_signal_3095), .B0_t (keyFF_outputPar[58]), .B0_f (new_AGEMA_signal_2534), .B1_t (new_AGEMA_signal_2535), .B1_f (new_AGEMA_signal_2536), .Z0_t (keyFF_inputPar[55]), .Z0_f (new_AGEMA_signal_3538), .Z1_t (new_AGEMA_signal_3539), .Z1_f (new_AGEMA_signal_3540) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[59]), .A0_f (new_AGEMA_signal_2543), .A1_t (new_AGEMA_signal_2544), .A1_f (new_AGEMA_signal_2545), .B0_t (key_s0_t[56]), .B0_f (key_s0_f[56]), .B1_t (key_s1_t[56]), .B1_f (key_s1_f[56]), .Z0_t (keyFF_MUX_inputPar_mux_inst_56_U1_X), .Z0_f (new_AGEMA_signal_2549), .Z1_t (new_AGEMA_signal_2550), .Z1_f (new_AGEMA_signal_2551) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_56_U1_X), .B0_f (new_AGEMA_signal_2549), .B1_t (new_AGEMA_signal_2550), .B1_f (new_AGEMA_signal_2551), .Z0_t (keyFF_MUX_inputPar_mux_inst_56_U1_Y), .Z0_f (new_AGEMA_signal_3096), .Z1_t (new_AGEMA_signal_3097), .Z1_f (new_AGEMA_signal_3098) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_56_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_56_U1_Y), .A0_f (new_AGEMA_signal_3096), .A1_t (new_AGEMA_signal_3097), .A1_f (new_AGEMA_signal_3098), .B0_t (keyFF_outputPar[59]), .B0_f (new_AGEMA_signal_2543), .B1_t (new_AGEMA_signal_2544), .B1_f (new_AGEMA_signal_2545), .Z0_t (keyFF_inputPar[56]), .Z0_f (new_AGEMA_signal_3541), .Z1_t (new_AGEMA_signal_3542), .Z1_f (new_AGEMA_signal_3543) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[60]), .A0_f (new_AGEMA_signal_2552), .A1_t (new_AGEMA_signal_2553), .A1_f (new_AGEMA_signal_2554), .B0_t (key_s0_t[57]), .B0_f (key_s0_f[57]), .B1_t (key_s1_t[57]), .B1_f (key_s1_f[57]), .Z0_t (keyFF_MUX_inputPar_mux_inst_57_U1_X), .Z0_f (new_AGEMA_signal_2558), .Z1_t (new_AGEMA_signal_2559), .Z1_f (new_AGEMA_signal_2560) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_57_U1_X), .B0_f (new_AGEMA_signal_2558), .B1_t (new_AGEMA_signal_2559), .B1_f (new_AGEMA_signal_2560), .Z0_t (keyFF_MUX_inputPar_mux_inst_57_U1_Y), .Z0_f (new_AGEMA_signal_3099), .Z1_t (new_AGEMA_signal_3100), .Z1_f (new_AGEMA_signal_3101) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_57_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_57_U1_Y), .A0_f (new_AGEMA_signal_3099), .A1_t (new_AGEMA_signal_3100), .A1_f (new_AGEMA_signal_3101), .B0_t (keyFF_outputPar[60]), .B0_f (new_AGEMA_signal_2552), .B1_t (new_AGEMA_signal_2553), .B1_f (new_AGEMA_signal_2554), .Z0_t (keyFF_inputPar[57]), .Z0_f (new_AGEMA_signal_3544), .Z1_t (new_AGEMA_signal_3545), .Z1_f (new_AGEMA_signal_3546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[61]), .A0_f (new_AGEMA_signal_2561), .A1_t (new_AGEMA_signal_2562), .A1_f (new_AGEMA_signal_2563), .B0_t (key_s0_t[58]), .B0_f (key_s0_f[58]), .B1_t (key_s1_t[58]), .B1_f (key_s1_f[58]), .Z0_t (keyFF_MUX_inputPar_mux_inst_58_U1_X), .Z0_f (new_AGEMA_signal_2567), .Z1_t (new_AGEMA_signal_2568), .Z1_f (new_AGEMA_signal_2569) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_58_U1_X), .B0_f (new_AGEMA_signal_2567), .B1_t (new_AGEMA_signal_2568), .B1_f (new_AGEMA_signal_2569), .Z0_t (keyFF_MUX_inputPar_mux_inst_58_U1_Y), .Z0_f (new_AGEMA_signal_3102), .Z1_t (new_AGEMA_signal_3103), .Z1_f (new_AGEMA_signal_3104) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_58_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_58_U1_Y), .A0_f (new_AGEMA_signal_3102), .A1_t (new_AGEMA_signal_3103), .A1_f (new_AGEMA_signal_3104), .B0_t (keyFF_outputPar[61]), .B0_f (new_AGEMA_signal_2561), .B1_t (new_AGEMA_signal_2562), .B1_f (new_AGEMA_signal_2563), .Z0_t (keyFF_inputPar[58]), .Z0_f (new_AGEMA_signal_3547), .Z1_t (new_AGEMA_signal_3548), .Z1_f (new_AGEMA_signal_3549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[62]), .A0_f (new_AGEMA_signal_2570), .A1_t (new_AGEMA_signal_2571), .A1_f (new_AGEMA_signal_2572), .B0_t (key_s0_t[59]), .B0_f (key_s0_f[59]), .B1_t (key_s1_t[59]), .B1_f (key_s1_f[59]), .Z0_t (keyFF_MUX_inputPar_mux_inst_59_U1_X), .Z0_f (new_AGEMA_signal_2576), .Z1_t (new_AGEMA_signal_2577), .Z1_f (new_AGEMA_signal_2578) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_59_U1_X), .B0_f (new_AGEMA_signal_2576), .B1_t (new_AGEMA_signal_2577), .B1_f (new_AGEMA_signal_2578), .Z0_t (keyFF_MUX_inputPar_mux_inst_59_U1_Y), .Z0_f (new_AGEMA_signal_3105), .Z1_t (new_AGEMA_signal_3106), .Z1_f (new_AGEMA_signal_3107) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_59_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_59_U1_Y), .A0_f (new_AGEMA_signal_3105), .A1_t (new_AGEMA_signal_3106), .A1_f (new_AGEMA_signal_3107), .B0_t (keyFF_outputPar[62]), .B0_f (new_AGEMA_signal_2570), .B1_t (new_AGEMA_signal_2571), .B1_f (new_AGEMA_signal_2572), .Z0_t (keyFF_inputPar[59]), .Z0_f (new_AGEMA_signal_3550), .Z1_t (new_AGEMA_signal_3551), .Z1_f (new_AGEMA_signal_3552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[63]), .A0_f (new_AGEMA_signal_2579), .A1_t (new_AGEMA_signal_2580), .A1_f (new_AGEMA_signal_2581), .B0_t (key_s0_t[60]), .B0_f (key_s0_f[60]), .B1_t (key_s1_t[60]), .B1_f (key_s1_f[60]), .Z0_t (keyFF_MUX_inputPar_mux_inst_60_U1_X), .Z0_f (new_AGEMA_signal_2585), .Z1_t (new_AGEMA_signal_2586), .Z1_f (new_AGEMA_signal_2587) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_60_U1_X), .B0_f (new_AGEMA_signal_2585), .B1_t (new_AGEMA_signal_2586), .B1_f (new_AGEMA_signal_2587), .Z0_t (keyFF_MUX_inputPar_mux_inst_60_U1_Y), .Z0_f (new_AGEMA_signal_3108), .Z1_t (new_AGEMA_signal_3109), .Z1_f (new_AGEMA_signal_3110) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_60_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_60_U1_Y), .A0_f (new_AGEMA_signal_3108), .A1_t (new_AGEMA_signal_3109), .A1_f (new_AGEMA_signal_3110), .B0_t (keyFF_outputPar[63]), .B0_f (new_AGEMA_signal_2579), .B1_t (new_AGEMA_signal_2580), .B1_f (new_AGEMA_signal_2581), .Z0_t (keyFF_inputPar[60]), .Z0_f (new_AGEMA_signal_3553), .Z1_t (new_AGEMA_signal_3554), .Z1_f (new_AGEMA_signal_3555) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[64]), .A0_f (new_AGEMA_signal_2588), .A1_t (new_AGEMA_signal_2589), .A1_f (new_AGEMA_signal_2590), .B0_t (key_s0_t[61]), .B0_f (key_s0_f[61]), .B1_t (key_s1_t[61]), .B1_f (key_s1_f[61]), .Z0_t (keyFF_MUX_inputPar_mux_inst_61_U1_X), .Z0_f (new_AGEMA_signal_2594), .Z1_t (new_AGEMA_signal_2595), .Z1_f (new_AGEMA_signal_2596) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_61_U1_X), .B0_f (new_AGEMA_signal_2594), .B1_t (new_AGEMA_signal_2595), .B1_f (new_AGEMA_signal_2596), .Z0_t (keyFF_MUX_inputPar_mux_inst_61_U1_Y), .Z0_f (new_AGEMA_signal_3111), .Z1_t (new_AGEMA_signal_3112), .Z1_f (new_AGEMA_signal_3113) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_61_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_61_U1_Y), .A0_f (new_AGEMA_signal_3111), .A1_t (new_AGEMA_signal_3112), .A1_f (new_AGEMA_signal_3113), .B0_t (keyFF_outputPar[64]), .B0_f (new_AGEMA_signal_2588), .B1_t (new_AGEMA_signal_2589), .B1_f (new_AGEMA_signal_2590), .Z0_t (keyFF_inputPar[61]), .Z0_f (new_AGEMA_signal_3556), .Z1_t (new_AGEMA_signal_3557), .Z1_f (new_AGEMA_signal_3558) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[65]), .A0_f (new_AGEMA_signal_2597), .A1_t (new_AGEMA_signal_2598), .A1_f (new_AGEMA_signal_2599), .B0_t (key_s0_t[62]), .B0_f (key_s0_f[62]), .B1_t (key_s1_t[62]), .B1_f (key_s1_f[62]), .Z0_t (keyFF_MUX_inputPar_mux_inst_62_U1_X), .Z0_f (new_AGEMA_signal_2603), .Z1_t (new_AGEMA_signal_2604), .Z1_f (new_AGEMA_signal_2605) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_62_U1_X), .B0_f (new_AGEMA_signal_2603), .B1_t (new_AGEMA_signal_2604), .B1_f (new_AGEMA_signal_2605), .Z0_t (keyFF_MUX_inputPar_mux_inst_62_U1_Y), .Z0_f (new_AGEMA_signal_3114), .Z1_t (new_AGEMA_signal_3115), .Z1_f (new_AGEMA_signal_3116) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_62_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_62_U1_Y), .A0_f (new_AGEMA_signal_3114), .A1_t (new_AGEMA_signal_3115), .A1_f (new_AGEMA_signal_3116), .B0_t (keyFF_outputPar[65]), .B0_f (new_AGEMA_signal_2597), .B1_t (new_AGEMA_signal_2598), .B1_f (new_AGEMA_signal_2599), .Z0_t (keyFF_inputPar[62]), .Z0_f (new_AGEMA_signal_3559), .Z1_t (new_AGEMA_signal_3560), .Z1_f (new_AGEMA_signal_3561) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[66]), .A0_f (new_AGEMA_signal_2606), .A1_t (new_AGEMA_signal_2607), .A1_f (new_AGEMA_signal_2608), .B0_t (key_s0_t[63]), .B0_f (key_s0_f[63]), .B1_t (key_s1_t[63]), .B1_f (key_s1_f[63]), .Z0_t (keyFF_MUX_inputPar_mux_inst_63_U1_X), .Z0_f (new_AGEMA_signal_2612), .Z1_t (new_AGEMA_signal_2613), .Z1_f (new_AGEMA_signal_2614) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_63_U1_X), .B0_f (new_AGEMA_signal_2612), .B1_t (new_AGEMA_signal_2613), .B1_f (new_AGEMA_signal_2614), .Z0_t (keyFF_MUX_inputPar_mux_inst_63_U1_Y), .Z0_f (new_AGEMA_signal_3117), .Z1_t (new_AGEMA_signal_3118), .Z1_f (new_AGEMA_signal_3119) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_63_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_63_U1_Y), .A0_f (new_AGEMA_signal_3117), .A1_t (new_AGEMA_signal_3118), .A1_f (new_AGEMA_signal_3119), .B0_t (keyFF_outputPar[66]), .B0_f (new_AGEMA_signal_2606), .B1_t (new_AGEMA_signal_2607), .B1_f (new_AGEMA_signal_2608), .Z0_t (keyFF_inputPar[63]), .Z0_f (new_AGEMA_signal_3562), .Z1_t (new_AGEMA_signal_3563), .Z1_f (new_AGEMA_signal_3564) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[67]), .A0_f (new_AGEMA_signal_2615), .A1_t (new_AGEMA_signal_2616), .A1_f (new_AGEMA_signal_2617), .B0_t (key_s0_t[64]), .B0_f (key_s0_f[64]), .B1_t (key_s1_t[64]), .B1_f (key_s1_f[64]), .Z0_t (keyFF_MUX_inputPar_mux_inst_64_U1_X), .Z0_f (new_AGEMA_signal_2621), .Z1_t (new_AGEMA_signal_2622), .Z1_f (new_AGEMA_signal_2623) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_64_U1_X), .B0_f (new_AGEMA_signal_2621), .B1_t (new_AGEMA_signal_2622), .B1_f (new_AGEMA_signal_2623), .Z0_t (keyFF_MUX_inputPar_mux_inst_64_U1_Y), .Z0_f (new_AGEMA_signal_3120), .Z1_t (new_AGEMA_signal_3121), .Z1_f (new_AGEMA_signal_3122) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_64_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_64_U1_Y), .A0_f (new_AGEMA_signal_3120), .A1_t (new_AGEMA_signal_3121), .A1_f (new_AGEMA_signal_3122), .B0_t (keyFF_outputPar[67]), .B0_f (new_AGEMA_signal_2615), .B1_t (new_AGEMA_signal_2616), .B1_f (new_AGEMA_signal_2617), .Z0_t (keyFF_inputPar[64]), .Z0_f (new_AGEMA_signal_3565), .Z1_t (new_AGEMA_signal_3566), .Z1_f (new_AGEMA_signal_3567) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[68]), .A0_f (new_AGEMA_signal_2624), .A1_t (new_AGEMA_signal_2625), .A1_f (new_AGEMA_signal_2626), .B0_t (key_s0_t[65]), .B0_f (key_s0_f[65]), .B1_t (key_s1_t[65]), .B1_f (key_s1_f[65]), .Z0_t (keyFF_MUX_inputPar_mux_inst_65_U1_X), .Z0_f (new_AGEMA_signal_2630), .Z1_t (new_AGEMA_signal_2631), .Z1_f (new_AGEMA_signal_2632) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_65_U1_X), .B0_f (new_AGEMA_signal_2630), .B1_t (new_AGEMA_signal_2631), .B1_f (new_AGEMA_signal_2632), .Z0_t (keyFF_MUX_inputPar_mux_inst_65_U1_Y), .Z0_f (new_AGEMA_signal_3123), .Z1_t (new_AGEMA_signal_3124), .Z1_f (new_AGEMA_signal_3125) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_65_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_65_U1_Y), .A0_f (new_AGEMA_signal_3123), .A1_t (new_AGEMA_signal_3124), .A1_f (new_AGEMA_signal_3125), .B0_t (keyFF_outputPar[68]), .B0_f (new_AGEMA_signal_2624), .B1_t (new_AGEMA_signal_2625), .B1_f (new_AGEMA_signal_2626), .Z0_t (keyFF_inputPar[65]), .Z0_f (new_AGEMA_signal_3568), .Z1_t (new_AGEMA_signal_3569), .Z1_f (new_AGEMA_signal_3570) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[69]), .A0_f (new_AGEMA_signal_2633), .A1_t (new_AGEMA_signal_2634), .A1_f (new_AGEMA_signal_2635), .B0_t (key_s0_t[66]), .B0_f (key_s0_f[66]), .B1_t (key_s1_t[66]), .B1_f (key_s1_f[66]), .Z0_t (keyFF_MUX_inputPar_mux_inst_66_U1_X), .Z0_f (new_AGEMA_signal_2639), .Z1_t (new_AGEMA_signal_2640), .Z1_f (new_AGEMA_signal_2641) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_66_U1_X), .B0_f (new_AGEMA_signal_2639), .B1_t (new_AGEMA_signal_2640), .B1_f (new_AGEMA_signal_2641), .Z0_t (keyFF_MUX_inputPar_mux_inst_66_U1_Y), .Z0_f (new_AGEMA_signal_3126), .Z1_t (new_AGEMA_signal_3127), .Z1_f (new_AGEMA_signal_3128) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_66_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_66_U1_Y), .A0_f (new_AGEMA_signal_3126), .A1_t (new_AGEMA_signal_3127), .A1_f (new_AGEMA_signal_3128), .B0_t (keyFF_outputPar[69]), .B0_f (new_AGEMA_signal_2633), .B1_t (new_AGEMA_signal_2634), .B1_f (new_AGEMA_signal_2635), .Z0_t (keyFF_inputPar[66]), .Z0_f (new_AGEMA_signal_3571), .Z1_t (new_AGEMA_signal_3572), .Z1_f (new_AGEMA_signal_3573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[70]), .A0_f (new_AGEMA_signal_2642), .A1_t (new_AGEMA_signal_2643), .A1_f (new_AGEMA_signal_2644), .B0_t (key_s0_t[67]), .B0_f (key_s0_f[67]), .B1_t (key_s1_t[67]), .B1_f (key_s1_f[67]), .Z0_t (keyFF_MUX_inputPar_mux_inst_67_U1_X), .Z0_f (new_AGEMA_signal_2648), .Z1_t (new_AGEMA_signal_2649), .Z1_f (new_AGEMA_signal_2650) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_67_U1_X), .B0_f (new_AGEMA_signal_2648), .B1_t (new_AGEMA_signal_2649), .B1_f (new_AGEMA_signal_2650), .Z0_t (keyFF_MUX_inputPar_mux_inst_67_U1_Y), .Z0_f (new_AGEMA_signal_3129), .Z1_t (new_AGEMA_signal_3130), .Z1_f (new_AGEMA_signal_3131) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_67_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_67_U1_Y), .A0_f (new_AGEMA_signal_3129), .A1_t (new_AGEMA_signal_3130), .A1_f (new_AGEMA_signal_3131), .B0_t (keyFF_outputPar[70]), .B0_f (new_AGEMA_signal_2642), .B1_t (new_AGEMA_signal_2643), .B1_f (new_AGEMA_signal_2644), .Z0_t (keyFF_inputPar[67]), .Z0_f (new_AGEMA_signal_3574), .Z1_t (new_AGEMA_signal_3575), .Z1_f (new_AGEMA_signal_3576) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[71]), .A0_f (new_AGEMA_signal_2651), .A1_t (new_AGEMA_signal_2652), .A1_f (new_AGEMA_signal_2653), .B0_t (key_s0_t[68]), .B0_f (key_s0_f[68]), .B1_t (key_s1_t[68]), .B1_f (key_s1_f[68]), .Z0_t (keyFF_MUX_inputPar_mux_inst_68_U1_X), .Z0_f (new_AGEMA_signal_2657), .Z1_t (new_AGEMA_signal_2658), .Z1_f (new_AGEMA_signal_2659) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_68_U1_X), .B0_f (new_AGEMA_signal_2657), .B1_t (new_AGEMA_signal_2658), .B1_f (new_AGEMA_signal_2659), .Z0_t (keyFF_MUX_inputPar_mux_inst_68_U1_Y), .Z0_f (new_AGEMA_signal_3132), .Z1_t (new_AGEMA_signal_3133), .Z1_f (new_AGEMA_signal_3134) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_68_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_68_U1_Y), .A0_f (new_AGEMA_signal_3132), .A1_t (new_AGEMA_signal_3133), .A1_f (new_AGEMA_signal_3134), .B0_t (keyFF_outputPar[71]), .B0_f (new_AGEMA_signal_2651), .B1_t (new_AGEMA_signal_2652), .B1_f (new_AGEMA_signal_2653), .Z0_t (keyFF_inputPar[68]), .Z0_f (new_AGEMA_signal_3577), .Z1_t (new_AGEMA_signal_3578), .Z1_f (new_AGEMA_signal_3579) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[72]), .A0_f (new_AGEMA_signal_2660), .A1_t (new_AGEMA_signal_2661), .A1_f (new_AGEMA_signal_2662), .B0_t (key_s0_t[69]), .B0_f (key_s0_f[69]), .B1_t (key_s1_t[69]), .B1_f (key_s1_f[69]), .Z0_t (keyFF_MUX_inputPar_mux_inst_69_U1_X), .Z0_f (new_AGEMA_signal_2666), .Z1_t (new_AGEMA_signal_2667), .Z1_f (new_AGEMA_signal_2668) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_69_U1_X), .B0_f (new_AGEMA_signal_2666), .B1_t (new_AGEMA_signal_2667), .B1_f (new_AGEMA_signal_2668), .Z0_t (keyFF_MUX_inputPar_mux_inst_69_U1_Y), .Z0_f (new_AGEMA_signal_3135), .Z1_t (new_AGEMA_signal_3136), .Z1_f (new_AGEMA_signal_3137) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_69_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_69_U1_Y), .A0_f (new_AGEMA_signal_3135), .A1_t (new_AGEMA_signal_3136), .A1_f (new_AGEMA_signal_3137), .B0_t (keyFF_outputPar[72]), .B0_f (new_AGEMA_signal_2660), .B1_t (new_AGEMA_signal_2661), .B1_f (new_AGEMA_signal_2662), .Z0_t (keyFF_inputPar[69]), .Z0_f (new_AGEMA_signal_3580), .Z1_t (new_AGEMA_signal_3581), .Z1_f (new_AGEMA_signal_3582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[73]), .A0_f (new_AGEMA_signal_2669), .A1_t (new_AGEMA_signal_2670), .A1_f (new_AGEMA_signal_2671), .B0_t (key_s0_t[70]), .B0_f (key_s0_f[70]), .B1_t (key_s1_t[70]), .B1_f (key_s1_f[70]), .Z0_t (keyFF_MUX_inputPar_mux_inst_70_U1_X), .Z0_f (new_AGEMA_signal_2675), .Z1_t (new_AGEMA_signal_2676), .Z1_f (new_AGEMA_signal_2677) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_70_U1_X), .B0_f (new_AGEMA_signal_2675), .B1_t (new_AGEMA_signal_2676), .B1_f (new_AGEMA_signal_2677), .Z0_t (keyFF_MUX_inputPar_mux_inst_70_U1_Y), .Z0_f (new_AGEMA_signal_3138), .Z1_t (new_AGEMA_signal_3139), .Z1_f (new_AGEMA_signal_3140) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_70_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_70_U1_Y), .A0_f (new_AGEMA_signal_3138), .A1_t (new_AGEMA_signal_3139), .A1_f (new_AGEMA_signal_3140), .B0_t (keyFF_outputPar[73]), .B0_f (new_AGEMA_signal_2669), .B1_t (new_AGEMA_signal_2670), .B1_f (new_AGEMA_signal_2671), .Z0_t (keyFF_inputPar[70]), .Z0_f (new_AGEMA_signal_3583), .Z1_t (new_AGEMA_signal_3584), .Z1_f (new_AGEMA_signal_3585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[74]), .A0_f (new_AGEMA_signal_2678), .A1_t (new_AGEMA_signal_2679), .A1_f (new_AGEMA_signal_2680), .B0_t (key_s0_t[71]), .B0_f (key_s0_f[71]), .B1_t (key_s1_t[71]), .B1_f (key_s1_f[71]), .Z0_t (keyFF_MUX_inputPar_mux_inst_71_U1_X), .Z0_f (new_AGEMA_signal_2684), .Z1_t (new_AGEMA_signal_2685), .Z1_f (new_AGEMA_signal_2686) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_71_U1_X), .B0_f (new_AGEMA_signal_2684), .B1_t (new_AGEMA_signal_2685), .B1_f (new_AGEMA_signal_2686), .Z0_t (keyFF_MUX_inputPar_mux_inst_71_U1_Y), .Z0_f (new_AGEMA_signal_3141), .Z1_t (new_AGEMA_signal_3142), .Z1_f (new_AGEMA_signal_3143) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_71_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_71_U1_Y), .A0_f (new_AGEMA_signal_3141), .A1_t (new_AGEMA_signal_3142), .A1_f (new_AGEMA_signal_3143), .B0_t (keyFF_outputPar[74]), .B0_f (new_AGEMA_signal_2678), .B1_t (new_AGEMA_signal_2679), .B1_f (new_AGEMA_signal_2680), .Z0_t (keyFF_inputPar[71]), .Z0_f (new_AGEMA_signal_3586), .Z1_t (new_AGEMA_signal_3587), .Z1_f (new_AGEMA_signal_3588) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_XOR1_U1 ( .A0_t (keyFF_outputPar[75]), .A0_f (new_AGEMA_signal_2687), .A1_t (new_AGEMA_signal_2688), .A1_f (new_AGEMA_signal_2689), .B0_t (key_s0_t[72]), .B0_f (key_s0_f[72]), .B1_t (key_s1_t[72]), .B1_f (key_s1_f[72]), .Z0_t (keyFF_MUX_inputPar_mux_inst_72_U1_X), .Z0_f (new_AGEMA_signal_2693), .Z1_t (new_AGEMA_signal_2694), .Z1_f (new_AGEMA_signal_2695) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_72_U1_X), .B0_f (new_AGEMA_signal_2693), .B1_t (new_AGEMA_signal_2694), .B1_f (new_AGEMA_signal_2695), .Z0_t (keyFF_MUX_inputPar_mux_inst_72_U1_Y), .Z0_f (new_AGEMA_signal_3144), .Z1_t (new_AGEMA_signal_3145), .Z1_f (new_AGEMA_signal_3146) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_72_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_72_U1_Y), .A0_f (new_AGEMA_signal_3144), .A1_t (new_AGEMA_signal_3145), .A1_f (new_AGEMA_signal_3146), .B0_t (keyFF_outputPar[75]), .B0_f (new_AGEMA_signal_2687), .B1_t (new_AGEMA_signal_2688), .B1_f (new_AGEMA_signal_2689), .Z0_t (keyFF_inputPar[72]), .Z0_f (new_AGEMA_signal_3589), .Z1_t (new_AGEMA_signal_3590), .Z1_f (new_AGEMA_signal_3591) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_XOR1_U1 ( .A0_t (roundkey[0]), .A0_f (new_AGEMA_signal_1452), .A1_t (new_AGEMA_signal_1453), .A1_f (new_AGEMA_signal_1454), .B0_t (key_s0_t[73]), .B0_f (key_s0_f[73]), .B1_t (key_s1_t[73]), .B1_f (key_s1_f[73]), .Z0_t (keyFF_MUX_inputPar_mux_inst_73_U1_X), .Z0_f (new_AGEMA_signal_2699), .Z1_t (new_AGEMA_signal_2700), .Z1_f (new_AGEMA_signal_2701) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_73_U1_X), .B0_f (new_AGEMA_signal_2699), .B1_t (new_AGEMA_signal_2700), .B1_f (new_AGEMA_signal_2701), .Z0_t (keyFF_MUX_inputPar_mux_inst_73_U1_Y), .Z0_f (new_AGEMA_signal_3147), .Z1_t (new_AGEMA_signal_3148), .Z1_f (new_AGEMA_signal_3149) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_73_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_73_U1_Y), .A0_f (new_AGEMA_signal_3147), .A1_t (new_AGEMA_signal_3148), .A1_f (new_AGEMA_signal_3149), .B0_t (roundkey[0]), .B0_f (new_AGEMA_signal_1452), .B1_t (new_AGEMA_signal_1453), .B1_f (new_AGEMA_signal_1454), .Z0_t (keyFF_inputPar[73]), .Z0_f (new_AGEMA_signal_3592), .Z1_t (new_AGEMA_signal_3593), .Z1_f (new_AGEMA_signal_3594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_XOR1_U1 ( .A0_t (roundkey[1]), .A0_f (new_AGEMA_signal_1434), .A1_t (new_AGEMA_signal_1435), .A1_f (new_AGEMA_signal_1436), .B0_t (key_s0_t[74]), .B0_f (key_s0_f[74]), .B1_t (key_s1_t[74]), .B1_f (key_s1_f[74]), .Z0_t (keyFF_MUX_inputPar_mux_inst_74_U1_X), .Z0_f (new_AGEMA_signal_2705), .Z1_t (new_AGEMA_signal_2706), .Z1_f (new_AGEMA_signal_2707) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_74_U1_X), .B0_f (new_AGEMA_signal_2705), .B1_t (new_AGEMA_signal_2706), .B1_f (new_AGEMA_signal_2707), .Z0_t (keyFF_MUX_inputPar_mux_inst_74_U1_Y), .Z0_f (new_AGEMA_signal_3150), .Z1_t (new_AGEMA_signal_3151), .Z1_f (new_AGEMA_signal_3152) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_74_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_74_U1_Y), .A0_f (new_AGEMA_signal_3150), .A1_t (new_AGEMA_signal_3151), .A1_f (new_AGEMA_signal_3152), .B0_t (roundkey[1]), .B0_f (new_AGEMA_signal_1434), .B1_t (new_AGEMA_signal_1435), .B1_f (new_AGEMA_signal_1436), .Z0_t (keyFF_inputPar[74]), .Z0_f (new_AGEMA_signal_3595), .Z1_t (new_AGEMA_signal_3596), .Z1_f (new_AGEMA_signal_3597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_XOR1_U1 ( .A0_t (roundkey[2]), .A0_f (new_AGEMA_signal_1443), .A1_t (new_AGEMA_signal_1444), .A1_f (new_AGEMA_signal_1445), .B0_t (key_s0_t[75]), .B0_f (key_s0_f[75]), .B1_t (key_s1_t[75]), .B1_f (key_s1_f[75]), .Z0_t (keyFF_MUX_inputPar_mux_inst_75_U1_X), .Z0_f (new_AGEMA_signal_2711), .Z1_t (new_AGEMA_signal_2712), .Z1_f (new_AGEMA_signal_2713) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_75_U1_X), .B0_f (new_AGEMA_signal_2711), .B1_t (new_AGEMA_signal_2712), .B1_f (new_AGEMA_signal_2713), .Z0_t (keyFF_MUX_inputPar_mux_inst_75_U1_Y), .Z0_f (new_AGEMA_signal_3153), .Z1_t (new_AGEMA_signal_3154), .Z1_f (new_AGEMA_signal_3155) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_75_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_75_U1_Y), .A0_f (new_AGEMA_signal_3153), .A1_t (new_AGEMA_signal_3154), .A1_f (new_AGEMA_signal_3155), .B0_t (roundkey[2]), .B0_f (new_AGEMA_signal_1443), .B1_t (new_AGEMA_signal_1444), .B1_f (new_AGEMA_signal_1445), .Z0_t (keyFF_inputPar[75]), .Z0_f (new_AGEMA_signal_3598), .Z1_t (new_AGEMA_signal_3599), .Z1_f (new_AGEMA_signal_3600) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_XOR1_U1 ( .A0_t (sboxOut[0]), .A0_f (new_AGEMA_signal_4491), .A1_t (new_AGEMA_signal_4492), .A1_f (new_AGEMA_signal_4493), .B0_t (key_s0_t[76]), .B0_f (key_s0_f[76]), .B1_t (key_s1_t[76]), .B1_f (key_s1_f[76]), .Z0_t (keyFF_MUX_inputPar_mux_inst_76_U1_X), .Z0_f (new_AGEMA_signal_4499), .Z1_t (new_AGEMA_signal_4500), .Z1_f (new_AGEMA_signal_4501) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_76_U1_X), .B0_f (new_AGEMA_signal_4499), .B1_t (new_AGEMA_signal_4500), .B1_f (new_AGEMA_signal_4501), .Z0_t (keyFF_MUX_inputPar_mux_inst_76_U1_Y), .Z0_f (new_AGEMA_signal_4513), .Z1_t (new_AGEMA_signal_4514), .Z1_f (new_AGEMA_signal_4515) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_76_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_76_U1_Y), .A0_f (new_AGEMA_signal_4513), .A1_t (new_AGEMA_signal_4514), .A1_f (new_AGEMA_signal_4515), .B0_t (sboxOut[0]), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (keyFF_inputPar[76]), .Z0_f (new_AGEMA_signal_4526), .Z1_t (new_AGEMA_signal_4527), .Z1_f (new_AGEMA_signal_4528) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_XOR1_U1 ( .A0_t (sboxOut[1]), .A0_f (new_AGEMA_signal_4550), .A1_t (new_AGEMA_signal_4551), .A1_f (new_AGEMA_signal_4552), .B0_t (key_s0_t[77]), .B0_f (key_s0_f[77]), .B1_t (key_s1_t[77]), .B1_f (key_s1_f[77]), .Z0_t (keyFF_MUX_inputPar_mux_inst_77_U1_X), .Z0_f (new_AGEMA_signal_4562), .Z1_t (new_AGEMA_signal_4563), .Z1_f (new_AGEMA_signal_4564) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_77_U1_X), .B0_f (new_AGEMA_signal_4562), .B1_t (new_AGEMA_signal_4563), .B1_f (new_AGEMA_signal_4564), .Z0_t (keyFF_MUX_inputPar_mux_inst_77_U1_Y), .Z0_f (new_AGEMA_signal_4580), .Z1_t (new_AGEMA_signal_4581), .Z1_f (new_AGEMA_signal_4582) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_77_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_77_U1_Y), .A0_f (new_AGEMA_signal_4580), .A1_t (new_AGEMA_signal_4581), .A1_f (new_AGEMA_signal_4582), .B0_t (sboxOut[1]), .B0_f (new_AGEMA_signal_4550), .B1_t (new_AGEMA_signal_4551), .B1_f (new_AGEMA_signal_4552), .Z0_t (keyFF_inputPar[77]), .Z0_f (new_AGEMA_signal_4601), .Z1_t (new_AGEMA_signal_4602), .Z1_f (new_AGEMA_signal_4603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_XOR1_U1 ( .A0_t (sboxOut[2]), .A0_f (new_AGEMA_signal_4547), .A1_t (new_AGEMA_signal_4548), .A1_f (new_AGEMA_signal_4549), .B0_t (key_s0_t[78]), .B0_f (key_s0_f[78]), .B1_t (key_s1_t[78]), .B1_f (key_s1_f[78]), .Z0_t (keyFF_MUX_inputPar_mux_inst_78_U1_X), .Z0_f (new_AGEMA_signal_4568), .Z1_t (new_AGEMA_signal_4569), .Z1_f (new_AGEMA_signal_4570) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_78_U1_X), .B0_f (new_AGEMA_signal_4568), .B1_t (new_AGEMA_signal_4569), .B1_f (new_AGEMA_signal_4570), .Z0_t (keyFF_MUX_inputPar_mux_inst_78_U1_Y), .Z0_f (new_AGEMA_signal_4583), .Z1_t (new_AGEMA_signal_4584), .Z1_f (new_AGEMA_signal_4585) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_78_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_78_U1_Y), .A0_f (new_AGEMA_signal_4583), .A1_t (new_AGEMA_signal_4584), .A1_f (new_AGEMA_signal_4585), .B0_t (sboxOut[2]), .B0_f (new_AGEMA_signal_4547), .B1_t (new_AGEMA_signal_4548), .B1_f (new_AGEMA_signal_4549), .Z0_t (keyFF_inputPar[78]), .Z0_f (new_AGEMA_signal_4604), .Z1_t (new_AGEMA_signal_4605), .Z1_f (new_AGEMA_signal_4606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_XOR1_U1 ( .A0_t (sboxOut[3]), .A0_f (new_AGEMA_signal_4571), .A1_t (new_AGEMA_signal_4572), .A1_f (new_AGEMA_signal_4573), .B0_t (key_s0_t[79]), .B0_f (key_s0_f[79]), .B1_t (key_s1_t[79]), .B1_f (key_s1_f[79]), .Z0_t (keyFF_MUX_inputPar_mux_inst_79_U1_X), .Z0_f (new_AGEMA_signal_4589), .Z1_t (new_AGEMA_signal_4590), .Z1_f (new_AGEMA_signal_4591) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (reset_t), .A1_f (reset_f), .B0_t (keyFF_MUX_inputPar_mux_inst_79_U1_X), .B0_f (new_AGEMA_signal_4589), .B1_t (new_AGEMA_signal_4590), .B1_f (new_AGEMA_signal_4591), .Z0_t (keyFF_MUX_inputPar_mux_inst_79_U1_Y), .Z0_f (new_AGEMA_signal_4607), .Z1_t (new_AGEMA_signal_4608), .Z1_f (new_AGEMA_signal_4609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keyFF_MUX_inputPar_mux_inst_79_U1_XOR2_U1 ( .A0_t (keyFF_MUX_inputPar_mux_inst_79_U1_Y), .A0_f (new_AGEMA_signal_4607), .A1_t (new_AGEMA_signal_4608), .A1_f (new_AGEMA_signal_4609), .B0_t (sboxOut[3]), .B0_f (new_AGEMA_signal_4571), .B1_t (new_AGEMA_signal_4572), .B1_f (new_AGEMA_signal_4573), .Z0_t (keyFF_inputPar[79]), .Z0_f (new_AGEMA_signal_4631), .Z1_t (new_AGEMA_signal_4632), .Z1_f (new_AGEMA_signal_4633) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR1_U1 ( .A0_t (sboxIn[2]), .A0_f (new_AGEMA_signal_4031), .A1_t (new_AGEMA_signal_4032), .A1_f (new_AGEMA_signal_4033), .B0_t (sboxIn[1]), .B0_f (new_AGEMA_signal_4028), .B1_t (new_AGEMA_signal_4029), .B1_f (new_AGEMA_signal_4030), .Z0_t (sboxInst_L0), .Z0_f (new_AGEMA_signal_4447), .Z1_t (new_AGEMA_signal_4448), .Z1_f (new_AGEMA_signal_4449) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR2_U1 ( .A0_t (sboxIn[1]), .A0_f (new_AGEMA_signal_4028), .A1_t (new_AGEMA_signal_4029), .A1_f (new_AGEMA_signal_4030), .B0_t (sboxIn[0]), .B0_f (new_AGEMA_signal_4025), .B1_t (new_AGEMA_signal_4026), .B1_f (new_AGEMA_signal_4027), .Z0_t (sboxInst_L1), .Z0_f (new_AGEMA_signal_4450), .Z1_t (new_AGEMA_signal_4451), .Z1_f (new_AGEMA_signal_4452) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR3_U1 ( .A0_t (sboxInst_L1), .A0_f (new_AGEMA_signal_4450), .A1_t (new_AGEMA_signal_4451), .A1_f (new_AGEMA_signal_4452), .B0_t (sboxIn[3]), .B0_f (new_AGEMA_signal_4034), .B1_t (new_AGEMA_signal_4035), .B1_f (new_AGEMA_signal_4036), .Z0_t (sboxInst_L2), .Z0_f (new_AGEMA_signal_4479), .Z1_t (new_AGEMA_signal_4480), .Z1_f (new_AGEMA_signal_4481) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) sboxInst_XOR16_U1 ( .A0_t (sboxInst_T0), .A0_f (new_AGEMA_signal_4488), .A1_t (new_AGEMA_signal_4489), .A1_f (new_AGEMA_signal_4490), .B0_t (sboxInst_L2), .B0_f (new_AGEMA_signal_4479), .B1_t (new_AGEMA_signal_4480), .B1_f (new_AGEMA_signal_4481), .Z0_t (sboxInst_Q2), .Z0_f (new_AGEMA_signal_4502), .Z1_t (new_AGEMA_signal_4503), .Z1_f (new_AGEMA_signal_4504) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR4_U1 ( .A0_t (sboxIn[3]), .A0_f (new_AGEMA_signal_4034), .A1_t (new_AGEMA_signal_4035), .A1_f (new_AGEMA_signal_4036), .B0_t (sboxIn[0]), .B0_f (new_AGEMA_signal_4025), .B1_t (new_AGEMA_signal_4026), .B1_f (new_AGEMA_signal_4027), .Z0_t (sboxInst_L3), .Z0_f (new_AGEMA_signal_4453), .Z1_t (new_AGEMA_signal_4454), .Z1_f (new_AGEMA_signal_4455) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR5_U1 ( .A0_t (sboxInst_L3), .A0_f (new_AGEMA_signal_4453), .A1_t (new_AGEMA_signal_4454), .A1_f (new_AGEMA_signal_4455), .B0_t (sboxInst_L0), .B0_f (new_AGEMA_signal_4447), .B1_t (new_AGEMA_signal_4448), .B1_f (new_AGEMA_signal_4449), .Z0_t (sboxInst_Q3), .Z0_f (new_AGEMA_signal_4482), .Z1_t (new_AGEMA_signal_4483), .Z1_f (new_AGEMA_signal_4484) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR6_U1 ( .A0_t (sboxIn[3]), .A0_f (new_AGEMA_signal_4034), .A1_t (new_AGEMA_signal_4035), .A1_f (new_AGEMA_signal_4036), .B0_t (sboxIn[1]), .B0_f (new_AGEMA_signal_4028), .B1_t (new_AGEMA_signal_4029), .B1_f (new_AGEMA_signal_4030), .Z0_t (sboxInst_L4), .Z0_f (new_AGEMA_signal_4456), .Z1_t (new_AGEMA_signal_4457), .Z1_f (new_AGEMA_signal_4458) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR7_U1 ( .A0_t (sboxInst_T0), .A0_f (new_AGEMA_signal_4488), .A1_t (new_AGEMA_signal_4489), .A1_f (new_AGEMA_signal_4490), .B0_t (sboxInst_T2), .B0_f (new_AGEMA_signal_4459), .B1_t (new_AGEMA_signal_4460), .B1_f (new_AGEMA_signal_4461), .Z0_t (sboxInst_L5), .Z0_f (new_AGEMA_signal_4505), .Z1_t (new_AGEMA_signal_4506), .Z1_f (new_AGEMA_signal_4507) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) sboxInst_XOR8_U1 ( .A0_t (sboxInst_L4), .A0_f (new_AGEMA_signal_4456), .A1_t (new_AGEMA_signal_4457), .A1_f (new_AGEMA_signal_4458), .B0_t (sboxInst_L5), .B0_f (new_AGEMA_signal_4505), .B1_t (new_AGEMA_signal_4506), .B1_f (new_AGEMA_signal_4507), .Z0_t (sboxInst_Q6), .Z0_f (new_AGEMA_signal_4516), .Z1_t (new_AGEMA_signal_4517), .Z1_f (new_AGEMA_signal_4518) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR9_U1 ( .A0_t (sboxInst_L1), .A0_f (new_AGEMA_signal_4450), .A1_t (new_AGEMA_signal_4451), .A1_f (new_AGEMA_signal_4452), .B0_t (sboxIn[2]), .B0_f (new_AGEMA_signal_4031), .B1_t (new_AGEMA_signal_4032), .B1_f (new_AGEMA_signal_4033), .Z0_t (sboxInst_Q7), .Z0_f (new_AGEMA_signal_4485), .Z1_t (new_AGEMA_signal_4486), .Z1_f (new_AGEMA_signal_4487) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) sboxInst_AND1_U1 ( .A0_t (sboxInst_L0), .A0_f (new_AGEMA_signal_4447), .A1_t (new_AGEMA_signal_4448), .A1_f (new_AGEMA_signal_4449), .B0_t (sboxIn[3]), .B0_f (new_AGEMA_signal_4034), .B1_t (new_AGEMA_signal_4035), .B1_f (new_AGEMA_signal_4036), .Z0_t (sboxInst_T0), .Z0_f (new_AGEMA_signal_4488), .Z1_t (new_AGEMA_signal_4489), .Z1_f (new_AGEMA_signal_4490) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND2_U1 ( .A0_t (sboxInst_Q2), .A0_f (new_AGEMA_signal_4502), .A1_t (new_AGEMA_signal_4503), .A1_f (new_AGEMA_signal_4504), .B0_t (sboxInst_Q3), .B0_f (new_AGEMA_signal_4482), .B1_t (new_AGEMA_signal_4483), .B1_f (new_AGEMA_signal_4484), .Z0_t (sboxInst_T1), .Z0_f (new_AGEMA_signal_4519), .Z1_t (new_AGEMA_signal_4520), .Z1_f (new_AGEMA_signal_4521) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND3_U1 ( .A0_t (sboxIn[1]), .A0_f (new_AGEMA_signal_4028), .A1_t (new_AGEMA_signal_4029), .A1_f (new_AGEMA_signal_4030), .B0_t (sboxIn[2]), .B0_f (new_AGEMA_signal_4031), .B1_t (new_AGEMA_signal_4032), .B1_f (new_AGEMA_signal_4033), .Z0_t (sboxInst_T2), .Z0_f (new_AGEMA_signal_4459), .Z1_t (new_AGEMA_signal_4460), .Z1_f (new_AGEMA_signal_4461) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_AND4_U1 ( .A0_t (sboxInst_Q6), .A0_f (new_AGEMA_signal_4516), .A1_t (new_AGEMA_signal_4517), .A1_f (new_AGEMA_signal_4518), .B0_t (sboxInst_Q7), .B0_f (new_AGEMA_signal_4485), .B1_t (new_AGEMA_signal_4486), .B1_f (new_AGEMA_signal_4487), .Z0_t (sboxInst_T3), .Z0_f (new_AGEMA_signal_4529), .Z1_t (new_AGEMA_signal_4530), .Z1_f (new_AGEMA_signal_4531) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR10_U1 ( .A0_t (sboxInst_L5), .A0_f (new_AGEMA_signal_4505), .A1_t (new_AGEMA_signal_4506), .A1_f (new_AGEMA_signal_4507), .B0_t (sboxInst_T3), .B0_f (new_AGEMA_signal_4529), .B1_t (new_AGEMA_signal_4530), .B1_f (new_AGEMA_signal_4531), .Z0_t (sboxInst_L7), .Z0_f (new_AGEMA_signal_4544), .Z1_t (new_AGEMA_signal_4545), .Z1_f (new_AGEMA_signal_4546) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR11_U1 ( .A0_t (sboxIn[0]), .A0_f (new_AGEMA_signal_4025), .A1_t (new_AGEMA_signal_4026), .A1_f (new_AGEMA_signal_4027), .B0_t (sboxInst_L7), .B0_f (new_AGEMA_signal_4544), .B1_t (new_AGEMA_signal_4545), .B1_f (new_AGEMA_signal_4546), .Z0_t (sboxOut[3]), .Z0_f (new_AGEMA_signal_4571), .Z1_t (new_AGEMA_signal_4572), .Z1_f (new_AGEMA_signal_4573) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR12_U1 ( .A0_t (sboxInst_L5), .A0_f (new_AGEMA_signal_4505), .A1_t (new_AGEMA_signal_4506), .A1_f (new_AGEMA_signal_4507), .B0_t (sboxInst_T1), .B0_f (new_AGEMA_signal_4519), .B1_t (new_AGEMA_signal_4520), .B1_f (new_AGEMA_signal_4521), .Z0_t (sboxInst_L8), .Z0_f (new_AGEMA_signal_4532), .Z1_t (new_AGEMA_signal_4533), .Z1_f (new_AGEMA_signal_4534) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR13_U1 ( .A0_t (sboxInst_L1), .A0_f (new_AGEMA_signal_4450), .A1_t (new_AGEMA_signal_4451), .A1_f (new_AGEMA_signal_4452), .B0_t (sboxInst_L8), .B0_f (new_AGEMA_signal_4532), .B1_t (new_AGEMA_signal_4533), .B1_f (new_AGEMA_signal_4534), .Z0_t (sboxOut[2]), .Z0_f (new_AGEMA_signal_4547), .Z1_t (new_AGEMA_signal_4548), .Z1_f (new_AGEMA_signal_4549) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR14_U1 ( .A0_t (sboxInst_L4), .A0_f (new_AGEMA_signal_4456), .A1_t (new_AGEMA_signal_4457), .A1_f (new_AGEMA_signal_4458), .B0_t (sboxInst_T3), .B0_f (new_AGEMA_signal_4529), .B1_t (new_AGEMA_signal_4530), .B1_f (new_AGEMA_signal_4531), .Z0_t (sboxOut[1]), .Z0_f (new_AGEMA_signal_4550), .Z1_t (new_AGEMA_signal_4551), .Z1_f (new_AGEMA_signal_4552) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) sboxInst_XOR15_U1 ( .A0_t (sboxInst_L3), .A0_f (new_AGEMA_signal_4453), .A1_t (new_AGEMA_signal_4454), .A1_f (new_AGEMA_signal_4455), .B0_t (sboxInst_T2), .B0_f (new_AGEMA_signal_4459), .B1_t (new_AGEMA_signal_4460), .B1_f (new_AGEMA_signal_4461), .Z0_t (sboxOut[0]), .Z0_f (new_AGEMA_signal_4491), .Z1_t (new_AGEMA_signal_4492), .Z1_f (new_AGEMA_signal_4493) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_XOR1_U1 ( .A0_t (stateXORroundkey[0]), .A0_f (new_AGEMA_signal_1458), .A1_t (new_AGEMA_signal_1459), .A1_f (new_AGEMA_signal_1460), .B0_t (roundkey[3]), .B0_f (new_AGEMA_signal_1461), .B1_t (new_AGEMA_signal_1462), .B1_f (new_AGEMA_signal_1463), .Z0_t (MUX_sboxin_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_3156), .Z1_t (new_AGEMA_signal_3157), .Z1_f (new_AGEMA_signal_3158) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selSbox), .A1_f (new_AGEMA_signal_1487), .B0_t (MUX_sboxin_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_3156), .B1_t (new_AGEMA_signal_3157), .B1_f (new_AGEMA_signal_3158), .Z0_t (MUX_sboxin_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_3601), .Z1_t (new_AGEMA_signal_3602), .Z1_f (new_AGEMA_signal_3603) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_0_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_3601), .A1_t (new_AGEMA_signal_3602), .A1_f (new_AGEMA_signal_3603), .B0_t (stateXORroundkey[0]), .B0_f (new_AGEMA_signal_1458), .B1_t (new_AGEMA_signal_1459), .B1_f (new_AGEMA_signal_1460), .Z0_t (sboxIn[0]), .Z0_f (new_AGEMA_signal_4025), .Z1_t (new_AGEMA_signal_4026), .Z1_f (new_AGEMA_signal_4027) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_XOR1_U1 ( .A0_t (stateXORroundkey[1]), .A0_f (new_AGEMA_signal_1440), .A1_t (new_AGEMA_signal_1441), .A1_f (new_AGEMA_signal_1442), .B0_t (keyRegKS[1]), .B0_f (new_AGEMA_signal_3159), .B1_t (new_AGEMA_signal_3160), .B1_f (new_AGEMA_signal_3161), .Z0_t (MUX_sboxin_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_3162), .Z1_t (new_AGEMA_signal_3163), .Z1_f (new_AGEMA_signal_3164) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selSbox), .A1_f (new_AGEMA_signal_1487), .B0_t (MUX_sboxin_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_3162), .B1_t (new_AGEMA_signal_3163), .B1_f (new_AGEMA_signal_3164), .Z0_t (MUX_sboxin_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_3604), .Z1_t (new_AGEMA_signal_3605), .Z1_f (new_AGEMA_signal_3606) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_1_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_3604), .A1_t (new_AGEMA_signal_3605), .A1_f (new_AGEMA_signal_3606), .B0_t (stateXORroundkey[1]), .B0_f (new_AGEMA_signal_1440), .B1_t (new_AGEMA_signal_1441), .B1_f (new_AGEMA_signal_1442), .Z0_t (sboxIn[1]), .Z0_f (new_AGEMA_signal_4028), .Z1_t (new_AGEMA_signal_4029), .Z1_f (new_AGEMA_signal_4030) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_XOR1_U1 ( .A0_t (stateXORroundkey[2]), .A0_f (new_AGEMA_signal_1449), .A1_t (new_AGEMA_signal_1450), .A1_f (new_AGEMA_signal_1451), .B0_t (keyRegKS[2]), .B0_f (new_AGEMA_signal_3165), .B1_t (new_AGEMA_signal_3166), .B1_f (new_AGEMA_signal_3167), .Z0_t (MUX_sboxin_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_3168), .Z1_t (new_AGEMA_signal_3169), .Z1_f (new_AGEMA_signal_3170) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selSbox), .A1_f (new_AGEMA_signal_1487), .B0_t (MUX_sboxin_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_3168), .B1_t (new_AGEMA_signal_3169), .B1_f (new_AGEMA_signal_3170), .Z0_t (MUX_sboxin_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_3607), .Z1_t (new_AGEMA_signal_3608), .Z1_f (new_AGEMA_signal_3609) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_2_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_3607), .A1_t (new_AGEMA_signal_3608), .A1_f (new_AGEMA_signal_3609), .B0_t (stateXORroundkey[2]), .B0_f (new_AGEMA_signal_1449), .B1_t (new_AGEMA_signal_1450), .B1_f (new_AGEMA_signal_1451), .Z0_t (sboxIn[2]), .Z0_f (new_AGEMA_signal_4031), .Z1_t (new_AGEMA_signal_4032), .Z1_f (new_AGEMA_signal_4033) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_XOR1_U1 ( .A0_t (stateXORroundkey[3]), .A0_f (new_AGEMA_signal_1467), .A1_t (new_AGEMA_signal_1468), .A1_f (new_AGEMA_signal_1469), .B0_t (keyRegKS[3]), .B0_f (new_AGEMA_signal_3171), .B1_t (new_AGEMA_signal_3172), .B1_f (new_AGEMA_signal_3173), .Z0_t (MUX_sboxin_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_3174), .Z1_t (new_AGEMA_signal_3175), .Z1_f (new_AGEMA_signal_3176) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (selSbox), .A1_f (new_AGEMA_signal_1487), .B0_t (MUX_sboxin_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_3174), .B1_t (new_AGEMA_signal_3175), .B1_f (new_AGEMA_signal_3176), .Z0_t (MUX_sboxin_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_3610), .Z1_t (new_AGEMA_signal_3611), .Z1_f (new_AGEMA_signal_3612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_sboxin_mux_inst_3_U1_XOR2_U1 ( .A0_t (MUX_sboxin_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_3610), .A1_t (new_AGEMA_signal_3611), .A1_f (new_AGEMA_signal_3612), .B0_t (stateXORroundkey[3]), .B0_f (new_AGEMA_signal_1467), .B1_t (new_AGEMA_signal_1468), .B1_f (new_AGEMA_signal_1469), .Z0_t (sboxIn[3]), .Z0_f (new_AGEMA_signal_4034), .Z1_t (new_AGEMA_signal_4035), .Z1_f (new_AGEMA_signal_4036) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_XOR1_U1 ( .A0_t (sboxOut[0]), .A0_f (new_AGEMA_signal_4491), .A1_t (new_AGEMA_signal_4492), .A1_f (new_AGEMA_signal_4493), .B0_t (stateXORroundkey[0]), .B0_f (new_AGEMA_signal_1458), .B1_t (new_AGEMA_signal_1459), .B1_f (new_AGEMA_signal_1460), .Z0_t (MUX_serialIn_mux_inst_0_U1_X), .Z0_f (new_AGEMA_signal_4508), .Z1_t (new_AGEMA_signal_4509), .Z1_f (new_AGEMA_signal_4510) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intDone), .A1_f (new_AGEMA_signal_1480), .B0_t (MUX_serialIn_mux_inst_0_U1_X), .B0_f (new_AGEMA_signal_4508), .B1_t (new_AGEMA_signal_4509), .B1_f (new_AGEMA_signal_4510), .Z0_t (MUX_serialIn_mux_inst_0_U1_Y), .Z0_f (new_AGEMA_signal_4522), .Z1_t (new_AGEMA_signal_4523), .Z1_f (new_AGEMA_signal_4524) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_0_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_0_U1_Y), .A0_f (new_AGEMA_signal_4522), .A1_t (new_AGEMA_signal_4523), .A1_f (new_AGEMA_signal_4524), .B0_t (sboxOut[0]), .B0_f (new_AGEMA_signal_4491), .B1_t (new_AGEMA_signal_4492), .B1_f (new_AGEMA_signal_4493), .Z0_t (serialIn[0]), .Z0_f (new_AGEMA_signal_4535), .Z1_t (new_AGEMA_signal_4536), .Z1_f (new_AGEMA_signal_4537) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_XOR1_U1 ( .A0_t (sboxOut[1]), .A0_f (new_AGEMA_signal_4550), .A1_t (new_AGEMA_signal_4551), .A1_f (new_AGEMA_signal_4552), .B0_t (stateXORroundkey[1]), .B0_f (new_AGEMA_signal_1440), .B1_t (new_AGEMA_signal_1441), .B1_f (new_AGEMA_signal_1442), .Z0_t (MUX_serialIn_mux_inst_1_U1_X), .Z0_f (new_AGEMA_signal_4574), .Z1_t (new_AGEMA_signal_4575), .Z1_f (new_AGEMA_signal_4576) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intDone), .A1_f (new_AGEMA_signal_1480), .B0_t (MUX_serialIn_mux_inst_1_U1_X), .B0_f (new_AGEMA_signal_4574), .B1_t (new_AGEMA_signal_4575), .B1_f (new_AGEMA_signal_4576), .Z0_t (MUX_serialIn_mux_inst_1_U1_Y), .Z0_f (new_AGEMA_signal_4592), .Z1_t (new_AGEMA_signal_4593), .Z1_f (new_AGEMA_signal_4594) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_1_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_1_U1_Y), .A0_f (new_AGEMA_signal_4592), .A1_t (new_AGEMA_signal_4593), .A1_f (new_AGEMA_signal_4594), .B0_t (sboxOut[1]), .B0_f (new_AGEMA_signal_4550), .B1_t (new_AGEMA_signal_4551), .B1_f (new_AGEMA_signal_4552), .Z0_t (serialIn[1]), .Z0_f (new_AGEMA_signal_4610), .Z1_t (new_AGEMA_signal_4611), .Z1_f (new_AGEMA_signal_4612) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_XOR1_U1 ( .A0_t (sboxOut[2]), .A0_f (new_AGEMA_signal_4547), .A1_t (new_AGEMA_signal_4548), .A1_f (new_AGEMA_signal_4549), .B0_t (stateXORroundkey[2]), .B0_f (new_AGEMA_signal_1449), .B1_t (new_AGEMA_signal_1450), .B1_f (new_AGEMA_signal_1451), .Z0_t (MUX_serialIn_mux_inst_2_U1_X), .Z0_f (new_AGEMA_signal_4577), .Z1_t (new_AGEMA_signal_4578), .Z1_f (new_AGEMA_signal_4579) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intDone), .A1_f (new_AGEMA_signal_1480), .B0_t (MUX_serialIn_mux_inst_2_U1_X), .B0_f (new_AGEMA_signal_4577), .B1_t (new_AGEMA_signal_4578), .B1_f (new_AGEMA_signal_4579), .Z0_t (MUX_serialIn_mux_inst_2_U1_Y), .Z0_f (new_AGEMA_signal_4595), .Z1_t (new_AGEMA_signal_4596), .Z1_f (new_AGEMA_signal_4597) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_2_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_2_U1_Y), .A0_f (new_AGEMA_signal_4595), .A1_t (new_AGEMA_signal_4596), .A1_f (new_AGEMA_signal_4597), .B0_t (sboxOut[2]), .B0_f (new_AGEMA_signal_4547), .B1_t (new_AGEMA_signal_4548), .B1_f (new_AGEMA_signal_4549), .Z0_t (serialIn[2]), .Z0_f (new_AGEMA_signal_4613), .Z1_t (new_AGEMA_signal_4614), .Z1_f (new_AGEMA_signal_4615) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_XOR1_U1 ( .A0_t (sboxOut[3]), .A0_f (new_AGEMA_signal_4571), .A1_t (new_AGEMA_signal_4572), .A1_f (new_AGEMA_signal_4573), .B0_t (stateXORroundkey[3]), .B0_f (new_AGEMA_signal_1467), .B1_t (new_AGEMA_signal_1468), .B1_f (new_AGEMA_signal_1469), .Z0_t (MUX_serialIn_mux_inst_3_U1_X), .Z0_f (new_AGEMA_signal_4598), .Z1_t (new_AGEMA_signal_4599), .Z1_f (new_AGEMA_signal_4600) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_AND1_U1 ( .A0_t (1'b0), .A0_f (1'b1), .A1_t (intDone), .A1_f (new_AGEMA_signal_1480), .B0_t (MUX_serialIn_mux_inst_3_U1_X), .B0_f (new_AGEMA_signal_4598), .B1_t (new_AGEMA_signal_4599), .B1_f (new_AGEMA_signal_4600), .Z0_t (MUX_serialIn_mux_inst_3_U1_Y), .Z0_f (new_AGEMA_signal_4616), .Z1_t (new_AGEMA_signal_4617), .Z1_f (new_AGEMA_signal_4618) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) MUX_serialIn_mux_inst_3_U1_XOR2_U1 ( .A0_t (MUX_serialIn_mux_inst_3_U1_Y), .A0_f (new_AGEMA_signal_4616), .A1_t (new_AGEMA_signal_4617), .A1_f (new_AGEMA_signal_4618), .B0_t (sboxOut[3]), .B0_f (new_AGEMA_signal_4571), .B1_t (new_AGEMA_signal_4572), .B1_f (new_AGEMA_signal_4573), .Z0_t (serialIn[3]), .Z0_f (new_AGEMA_signal_4634), .Z1_t (new_AGEMA_signal_4635), .Z1_f (new_AGEMA_signal_4636) ) ;

    /* register cells */
endmodule
