/* modified netlist. Source: module Midori64 in file /mnt/c/Users/amirm/Desktop/Papers_in_progress/SAUBER/Design for our FPGA/13-Midori64_round_based_enc_dec_PortParallel/4-AGEMA/Midori64.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module Midori64_SAUBER_Pipeline_d1 (DataIn, key, reset, enc_dec, DataOut, done);
    input [63:0] DataIn ;
    input [127:0] key ;
    input reset ;
    input enc_dec ;
    output [63:0] DataOut ;
    output done ;
    wire controller_n2 ;
    wire controller_n1 ;
    wire controller_roundCounter_n15 ;
    wire controller_roundCounter_n14 ;
    wire controller_roundCounter_n13 ;
    wire controller_roundCounter_n8 ;
    wire controller_roundCounter_n4 ;
    wire controller_roundCounter_n5 ;
    wire controller_roundCounter_n6 ;
    wire controller_roundCounter_N7 ;
    wire controller_roundCounter_U9_Y ;
    wire controller_roundCounter_U9_X ;
    wire controller_roundCounter_U11_Y ;
    wire controller_roundCounter_U11_X ;
    wire controller_roundCounter_U15_Y ;
    wire controller_roundCounter_U15_X ;
    wire Midori_rounds_n16 ;
    wire Midori_rounds_n15 ;
    wire Midori_rounds_n14 ;
    wire Midori_rounds_n13 ;
    wire Midori_rounds_n12 ;
    wire Midori_rounds_n11 ;
    wire Midori_rounds_n10 ;
    wire Midori_rounds_n9 ;
    wire Midori_rounds_n8 ;
    wire Midori_rounds_n7 ;
    wire Midori_rounds_n6 ;
    wire Midori_rounds_n5 ;
    wire Midori_rounds_n4 ;
    wire Midori_rounds_n3 ;
    wire Midori_rounds_n2 ;
    wire Midori_rounds_n1 ;
    wire Midori_rounds_constant_MUX_n139 ;
    wire Midori_rounds_constant_MUX_n138 ;
    wire Midori_rounds_constant_MUX_n137 ;
    wire Midori_rounds_constant_MUX_n136 ;
    wire Midori_rounds_constant_MUX_n134 ;
    wire Midori_rounds_constant_MUX_n133 ;
    wire Midori_rounds_constant_MUX_n132 ;
    wire Midori_rounds_constant_MUX_n131 ;
    wire Midori_rounds_constant_MUX_n130 ;
    wire Midori_rounds_constant_MUX_n129 ;
    wire Midori_rounds_constant_MUX_n128 ;
    wire Midori_rounds_constant_MUX_n126 ;
    wire Midori_rounds_constant_MUX_n125 ;
    wire Midori_rounds_constant_MUX_n124 ;
    wire Midori_rounds_constant_MUX_n123 ;
    wire Midori_rounds_constant_MUX_n122 ;
    wire Midori_rounds_constant_MUX_n120 ;
    wire Midori_rounds_constant_MUX_n119 ;
    wire Midori_rounds_constant_MUX_n118 ;
    wire Midori_rounds_constant_MUX_n117 ;
    wire Midori_rounds_constant_MUX_n116 ;
    wire Midori_rounds_constant_MUX_n115 ;
    wire Midori_rounds_constant_MUX_n114 ;
    wire Midori_rounds_constant_MUX_n113 ;
    wire Midori_rounds_constant_MUX_n110 ;
    wire Midori_rounds_constant_MUX_n109 ;
    wire Midori_rounds_constant_MUX_n108 ;
    wire Midori_rounds_constant_MUX_n107 ;
    wire Midori_rounds_constant_MUX_n106 ;
    wire Midori_rounds_constant_MUX_n104 ;
    wire Midori_rounds_constant_MUX_n103 ;
    wire Midori_rounds_constant_MUX_n102 ;
    wire Midori_rounds_constant_MUX_n101 ;
    wire Midori_rounds_constant_MUX_n100 ;
    wire Midori_rounds_constant_MUX_n99 ;
    wire Midori_rounds_constant_MUX_n98 ;
    wire Midori_rounds_constant_MUX_n97 ;
    wire Midori_rounds_constant_MUX_n96 ;
    wire Midori_rounds_constant_MUX_n95 ;
    wire Midori_rounds_constant_MUX_n94 ;
    wire Midori_rounds_constant_MUX_n93 ;
    wire Midori_rounds_constant_MUX_n92 ;
    wire Midori_rounds_constant_MUX_n91 ;
    wire Midori_rounds_constant_MUX_n88 ;
    wire Midori_rounds_constant_MUX_n86 ;
    wire Midori_rounds_constant_MUX_n85 ;
    wire Midori_rounds_constant_MUX_n84 ;
    wire Midori_rounds_constant_MUX_n83 ;
    wire Midori_rounds_constant_MUX_n82 ;
    wire Midori_rounds_constant_MUX_n81 ;
    wire Midori_rounds_constant_MUX_n80 ;
    wire Midori_rounds_constant_MUX_n79 ;
    wire Midori_rounds_constant_MUX_n78 ;
    wire Midori_rounds_constant_MUX_n77 ;
    wire Midori_rounds_constant_MUX_n76 ;
    wire Midori_rounds_constant_MUX_n75 ;
    wire Midori_rounds_constant_MUX_n74 ;
    wire Midori_rounds_constant_MUX_n73 ;
    wire Midori_rounds_constant_MUX_n72 ;
    wire Midori_rounds_constant_MUX_n70 ;
    wire Midori_rounds_constant_MUX_n69 ;
    wire Midori_rounds_constant_MUX_n68 ;
    wire Midori_rounds_constant_MUX_n66 ;
    wire Midori_rounds_constant_MUX_n64 ;
    wire Midori_rounds_constant_MUX_n62 ;
    wire Midori_rounds_constant_MUX_n61 ;
    wire Midori_rounds_constant_MUX_n60 ;
    wire Midori_rounds_constant_MUX_n59 ;
    wire Midori_rounds_constant_MUX_n58 ;
    wire Midori_rounds_constant_MUX_n57 ;
    wire Midori_rounds_constant_MUX_n56 ;
    wire Midori_rounds_constant_MUX_n55 ;
    wire Midori_rounds_constant_MUX_n54 ;
    wire Midori_rounds_constant_MUX_n53 ;
    wire Midori_rounds_constant_MUX_n52 ;
    wire Midori_rounds_constant_MUX_n51 ;
    wire Midori_rounds_constant_MUX_n50 ;
    wire Midori_rounds_constant_MUX_n49 ;
    wire Midori_rounds_constant_MUX_n48 ;
    wire Midori_rounds_constant_MUX_n47 ;
    wire Midori_rounds_constant_MUX_n46 ;
    wire Midori_rounds_constant_MUX_n42 ;
    wire Midori_rounds_constant_MUX_n40 ;
    wire Midori_rounds_constant_MUX_n37 ;
    wire Midori_rounds_constant_MUX_n36 ;
    wire Midori_rounds_constant_MUX_n35 ;
    wire Midori_rounds_constant_MUX_n34 ;
    wire Midori_rounds_constant_MUX_n33 ;
    wire Midori_rounds_constant_MUX_n32 ;
    wire Midori_rounds_constant_MUX_n31 ;
    wire Midori_rounds_constant_MUX_n30 ;
    wire Midori_rounds_constant_MUX_n29 ;
    wire Midori_rounds_constant_MUX_n28 ;
    wire Midori_rounds_constant_MUX_n27 ;
    wire Midori_rounds_constant_MUX_n25 ;
    wire Midori_rounds_constant_MUX_n24 ;
    wire Midori_rounds_constant_MUX_n23 ;
    wire Midori_rounds_constant_MUX_n22 ;
    wire Midori_rounds_constant_MUX_n121 ;
    wire Midori_rounds_constant_MUX_n112 ;
    wire Midori_rounds_constant_MUX_n43 ;
    wire Midori_rounds_constant_MUX_n111 ;
    wire Midori_rounds_constant_MUX_U53_Y ;
    wire Midori_rounds_constant_MUX_U53_X ;
    wire Midori_rounds_constant_MUX_U119_Y ;
    wire Midori_rounds_constant_MUX_U119_X ;
    wire Midori_rounds_MUXInst_mux_inst_0_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_0_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_1_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_1_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_2_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_2_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_3_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_3_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_4_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_4_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_5_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_5_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_6_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_6_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_7_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_7_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_8_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_8_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_9_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_9_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_10_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_10_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_11_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_11_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_12_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_12_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_13_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_13_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_14_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_14_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_15_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_15_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_16_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_16_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_17_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_17_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_18_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_18_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_19_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_19_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_20_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_20_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_21_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_21_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_22_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_22_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_23_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_23_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_24_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_24_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_25_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_25_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_26_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_26_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_27_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_27_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_28_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_28_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_29_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_29_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_30_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_30_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_31_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_31_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_32_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_32_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_33_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_33_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_34_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_34_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_35_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_35_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_36_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_36_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_37_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_37_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_38_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_38_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_39_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_39_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_40_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_40_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_41_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_41_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_42_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_42_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_43_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_43_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_44_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_44_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_45_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_45_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_46_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_46_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_47_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_47_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_48_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_48_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_49_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_49_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_50_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_50_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_51_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_51_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_52_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_52_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_53_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_53_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_54_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_54_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_55_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_55_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_56_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_56_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_57_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_57_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_58_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_58_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_59_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_59_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_60_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_60_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_61_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_61_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_62_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_62_U1_X ;
    wire Midori_rounds_MUXInst_mux_inst_63_U1_Y ;
    wire Midori_rounds_MUXInst_mux_inst_63_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X ;
    wire Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y ;
    wire Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_0_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_1_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_2_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_3_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_4_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_5_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_6_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_7_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_8_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_9_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_10_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_11_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_12_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_13_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n12 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n6 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_14_n1 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n15 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n14 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n13 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n11 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n10 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n9 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n8 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n7 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n5 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n3 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n2 ;
    wire Midori_rounds_sub_sBox_PRINCE_15_n1 ;
    wire Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_0_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_1_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_2_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_3_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_4_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_5_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_6_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_7_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_8_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_9_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_10_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_11_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_12_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_13_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_14_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_15_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_16_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_17_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_18_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_19_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_20_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_21_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_22_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_23_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_24_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_25_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_26_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_27_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_28_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_29_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_30_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_31_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_32_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_33_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_34_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_35_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_36_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_37_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_38_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_39_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_40_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_41_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_42_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_43_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_44_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_45_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_46_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_47_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_48_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_49_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_50_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_51_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_52_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_53_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_54_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_55_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_56_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_57_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_58_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_59_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_60_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_61_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_62_U1_X ;
    wire Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y ;
    wire Midori_rounds_mul_input_Inst_mux_inst_63_U1_X ;
    wire Midori_rounds_mul_MC1_n8 ;
    wire Midori_rounds_mul_MC1_n7 ;
    wire Midori_rounds_mul_MC1_n6 ;
    wire Midori_rounds_mul_MC1_n5 ;
    wire Midori_rounds_mul_MC1_n4 ;
    wire Midori_rounds_mul_MC1_n3 ;
    wire Midori_rounds_mul_MC1_n2 ;
    wire Midori_rounds_mul_MC1_n1 ;
    wire Midori_rounds_mul_MC2_n8 ;
    wire Midori_rounds_mul_MC2_n7 ;
    wire Midori_rounds_mul_MC2_n6 ;
    wire Midori_rounds_mul_MC2_n5 ;
    wire Midori_rounds_mul_MC2_n4 ;
    wire Midori_rounds_mul_MC2_n3 ;
    wire Midori_rounds_mul_MC2_n2 ;
    wire Midori_rounds_mul_MC2_n1 ;
    wire Midori_rounds_mul_MC3_n8 ;
    wire Midori_rounds_mul_MC3_n7 ;
    wire Midori_rounds_mul_MC3_n6 ;
    wire Midori_rounds_mul_MC3_n5 ;
    wire Midori_rounds_mul_MC3_n4 ;
    wire Midori_rounds_mul_MC3_n3 ;
    wire Midori_rounds_mul_MC3_n2 ;
    wire Midori_rounds_mul_MC3_n1 ;
    wire Midori_rounds_mul_MC4_n8 ;
    wire Midori_rounds_mul_MC4_n7 ;
    wire Midori_rounds_mul_MC4_n6 ;
    wire Midori_rounds_mul_MC4_n5 ;
    wire Midori_rounds_mul_MC4_n4 ;
    wire Midori_rounds_mul_MC4_n3 ;
    wire Midori_rounds_mul_MC4_n2 ;
    wire Midori_rounds_mul_MC4_n1 ;
    wire Midori_rounds_Res_Inst_mux_inst_0_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_0_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_1_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_1_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_2_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_2_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_3_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_3_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_4_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_4_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_5_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_5_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_6_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_6_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_7_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_7_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_8_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_8_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_9_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_9_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_10_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_10_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_11_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_11_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_12_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_12_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_13_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_13_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_14_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_14_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_15_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_15_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_16_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_16_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_17_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_17_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_18_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_18_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_19_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_19_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_20_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_20_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_21_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_21_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_22_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_22_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_23_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_23_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_24_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_24_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_25_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_25_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_26_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_26_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_27_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_27_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_28_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_28_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_29_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_29_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_30_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_30_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_31_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_31_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_32_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_32_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_33_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_33_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_34_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_34_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_35_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_35_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_36_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_36_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_37_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_37_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_38_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_38_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_39_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_39_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_40_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_40_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_41_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_41_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_42_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_42_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_43_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_43_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_44_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_44_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_45_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_45_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_46_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_46_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_47_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_47_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_48_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_48_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_49_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_49_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_50_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_50_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_51_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_51_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_52_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_52_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_53_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_53_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_54_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_54_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_55_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_55_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_56_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_56_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_57_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_57_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_58_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_58_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_59_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_59_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_60_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_60_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_61_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_61_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_62_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_62_U1_X ;
    wire Midori_rounds_Res_Inst_mux_inst_63_U1_Y ;
    wire Midori_rounds_Res_Inst_mux_inst_63_U1_X ;
    wire [63:0] wk ;
    wire [3:0] round_Signal ;
    wire [63:0] Midori_add_Result_Start ;
    wire [63:0] Midori_rounds_mul_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Inv_Result ;
    wire [63:0] Midori_rounds_mul_input ;
    wire [63:0] Midori_rounds_sub_ResultXORkey ;
    wire [63:0] Midori_rounds_SR_Result ;
    wire [63:0] Midori_rounds_roundReg_out ;
    wire [63:0] Midori_rounds_round_Result ;
    wire [63:0] Midori_rounds_SelectedKey ;
    wire [15:0] Midori_rounds_round_Constant ;

    /* cells in depth 0 */
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U64 ( .A0_t (key[127]), .B0_t (key[63]), .Z0_t (wk[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U63 ( .A0_t (key[126]), .B0_t (key[62]), .Z0_t (wk[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U62 ( .A0_t (key[125]), .B0_t (key[61]), .Z0_t (wk[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U61 ( .A0_t (key[124]), .B0_t (key[60]), .Z0_t (wk[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U60 ( .A0_t (key[123]), .B0_t (key[59]), .Z0_t (wk[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U59 ( .A0_t (key[122]), .B0_t (key[58]), .Z0_t (wk[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U58 ( .A0_t (key[121]), .B0_t (key[57]), .Z0_t (wk[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U57 ( .A0_t (key[120]), .B0_t (key[56]), .Z0_t (wk[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U56 ( .A0_t (key[119]), .B0_t (key[55]), .Z0_t (wk[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U55 ( .A0_t (key[118]), .B0_t (key[54]), .Z0_t (wk[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U54 ( .A0_t (key[117]), .B0_t (key[53]), .Z0_t (wk[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U53 ( .A0_t (key[116]), .B0_t (key[52]), .Z0_t (wk[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U52 ( .A0_t (key[115]), .B0_t (key[51]), .Z0_t (wk[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U51 ( .A0_t (key[114]), .B0_t (key[50]), .Z0_t (wk[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U50 ( .A0_t (key[113]), .B0_t (key[49]), .Z0_t (wk[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U49 ( .A0_t (key[112]), .B0_t (key[48]), .Z0_t (wk[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U48 ( .A0_t (key[111]), .B0_t (key[47]), .Z0_t (wk[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U47 ( .A0_t (key[110]), .B0_t (key[46]), .Z0_t (wk[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U46 ( .A0_t (key[109]), .B0_t (key[45]), .Z0_t (wk[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U45 ( .A0_t (key[108]), .B0_t (key[44]), .Z0_t (wk[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U44 ( .A0_t (key[107]), .B0_t (key[43]), .Z0_t (wk[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U43 ( .A0_t (key[106]), .B0_t (key[42]), .Z0_t (wk[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U42 ( .A0_t (key[105]), .B0_t (key[41]), .Z0_t (wk[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U41 ( .A0_t (key[104]), .B0_t (key[40]), .Z0_t (wk[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U40 ( .A0_t (key[103]), .B0_t (key[39]), .Z0_t (wk[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U39 ( .A0_t (key[102]), .B0_t (key[38]), .Z0_t (wk[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U38 ( .A0_t (key[101]), .B0_t (key[37]), .Z0_t (wk[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U37 ( .A0_t (key[100]), .B0_t (key[36]), .Z0_t (wk[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U36 ( .A0_t (key[99]), .B0_t (key[35]), .Z0_t (wk[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U35 ( .A0_t (key[98]), .B0_t (key[34]), .Z0_t (wk[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U34 ( .A0_t (key[97]), .B0_t (key[33]), .Z0_t (wk[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U33 ( .A0_t (key[96]), .B0_t (key[32]), .Z0_t (wk[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U32 ( .A0_t (key[95]), .B0_t (key[31]), .Z0_t (wk[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U31 ( .A0_t (key[94]), .B0_t (key[30]), .Z0_t (wk[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U30 ( .A0_t (key[93]), .B0_t (key[29]), .Z0_t (wk[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U29 ( .A0_t (key[92]), .B0_t (key[28]), .Z0_t (wk[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U28 ( .A0_t (key[91]), .B0_t (key[27]), .Z0_t (wk[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U27 ( .A0_t (key[90]), .B0_t (key[26]), .Z0_t (wk[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U26 ( .A0_t (key[89]), .B0_t (key[25]), .Z0_t (wk[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U25 ( .A0_t (key[88]), .B0_t (key[24]), .Z0_t (wk[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U24 ( .A0_t (key[87]), .B0_t (key[23]), .Z0_t (wk[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U23 ( .A0_t (key[86]), .B0_t (key[22]), .Z0_t (wk[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U22 ( .A0_t (key[85]), .B0_t (key[21]), .Z0_t (wk[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U21 ( .A0_t (key[84]), .B0_t (key[20]), .Z0_t (wk[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U20 ( .A0_t (key[83]), .B0_t (key[19]), .Z0_t (wk[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U19 ( .A0_t (key[82]), .B0_t (key[18]), .Z0_t (wk[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U18 ( .A0_t (key[81]), .B0_t (key[17]), .Z0_t (wk[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U17 ( .A0_t (key[80]), .B0_t (key[16]), .Z0_t (wk[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U16 ( .A0_t (key[79]), .B0_t (key[15]), .Z0_t (wk[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U15 ( .A0_t (key[78]), .B0_t (key[14]), .Z0_t (wk[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U14 ( .A0_t (key[77]), .B0_t (key[13]), .Z0_t (wk[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U13 ( .A0_t (key[76]), .B0_t (key[12]), .Z0_t (wk[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U12 ( .A0_t (key[75]), .B0_t (key[11]), .Z0_t (wk[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U11 ( .A0_t (key[74]), .B0_t (key[10]), .Z0_t (wk[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U10 ( .A0_t (key[73]), .B0_t (key[9]), .Z0_t (wk[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U9 ( .A0_t (key[72]), .B0_t (key[8]), .Z0_t (wk[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U8 ( .A0_t (key[71]), .B0_t (key[7]), .Z0_t (wk[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U7 ( .A0_t (key[70]), .B0_t (key[6]), .Z0_t (wk[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U6 ( .A0_t (key[69]), .B0_t (key[5]), .Z0_t (wk[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U5 ( .A0_t (key[68]), .B0_t (key[4]), .Z0_t (wk[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U4 ( .A0_t (key[67]), .B0_t (key[3]), .Z0_t (wk[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U3 ( .A0_t (key[66]), .B0_t (key[2]), .Z0_t (wk[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U2 ( .A0_t (key[65]), .B0_t (key[1]), .Z0_t (wk[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) keys_U1 ( .A0_t (key[64]), .B0_t (key[0]), .Z0_t (wk[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_U3 ( .A0_t (controller_n2), .B0_t (controller_n1), .Z0_t (done) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_U2 ( .A0_t (round_Signal[1]), .B0_t (round_Signal[0]), .Z0_t (controller_n1) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_U1 ( .A0_t (round_Signal[3]), .B0_t (round_Signal[2]), .Z0_t (controller_n2) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U10 ( .A0_t (round_Signal[2]), .B0_t (controller_roundCounter_n15), .Z0_t (controller_roundCounter_n5) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U8 ( .A0_t (round_Signal[1]), .B0_t (controller_roundCounter_n6), .Z0_t (controller_roundCounter_n15) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U7 ( .A0_t (reset), .B0_t (round_Signal[0]), .Z0_t (controller_roundCounter_n6) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U6 ( .A0_t (controller_roundCounter_n14), .B0_t (controller_roundCounter_n13), .Z0_t (controller_roundCounter_n4) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U5 ( .A0_t (round_Signal[2]), .B0_t (reset), .Z0_t (controller_roundCounter_n13) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U3 ( .A0_t (controller_roundCounter_N7), .B0_t (controller_roundCounter_n8), .Z0_t (controller_roundCounter_n14) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U2 ( .A0_t (reset), .B0_t (round_Signal[1]), .Z0_t (controller_roundCounter_n8) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U1 ( .A0_t (reset), .B0_t (round_Signal[0]), .Z0_t (controller_roundCounter_N7) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U9_XOR1_U1 ( .A0_t (controller_roundCounter_n5), .B0_t (controller_roundCounter_n4), .Z0_t (controller_roundCounter_U9_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U9_AND1_U1 ( .A0_t (round_Signal[3]), .B0_t (controller_roundCounter_U9_X), .Z0_t (controller_roundCounter_U9_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U9_XOR2_U1 ( .A0_t (controller_roundCounter_U9_Y), .B0_t (controller_roundCounter_n5), .Z0_t (round_Signal[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U11_XOR1_U1 ( .A0_t (controller_roundCounter_n6), .B0_t (controller_roundCounter_N7), .Z0_t (controller_roundCounter_U11_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U11_AND1_U1 ( .A0_t (round_Signal[1]), .B0_t (controller_roundCounter_U11_X), .Z0_t (controller_roundCounter_U11_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U11_XOR2_U1 ( .A0_t (controller_roundCounter_U11_Y), .B0_t (controller_roundCounter_n6), .Z0_t (round_Signal[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) controller_roundCounter_U15_XOR1_U1 ( .A0_t (controller_roundCounter_n14), .B0_t (controller_roundCounter_n15), .Z0_t (controller_roundCounter_U15_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) controller_roundCounter_U15_AND1_U1 ( .A0_t (round_Signal[2]), .B0_t (controller_roundCounter_U15_X), .Z0_t (controller_roundCounter_U15_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) controller_roundCounter_U15_XOR2_U1 ( .A0_t (controller_roundCounter_U15_Y), .B0_t (controller_roundCounter_n14), .Z0_t (round_Signal[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U128 ( .A0_t (wk[63]), .B0_t (DataIn[63]), .Z0_t (Midori_add_Result_Start[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U127 ( .A0_t (wk[62]), .B0_t (DataIn[62]), .Z0_t (Midori_add_Result_Start[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U126 ( .A0_t (wk[61]), .B0_t (DataIn[61]), .Z0_t (Midori_add_Result_Start[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U125 ( .A0_t (wk[60]), .B0_t (DataIn[60]), .Z0_t (Midori_add_Result_Start[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U124 ( .A0_t (wk[59]), .B0_t (DataIn[59]), .Z0_t (Midori_add_Result_Start[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U123 ( .A0_t (wk[58]), .B0_t (DataIn[58]), .Z0_t (Midori_add_Result_Start[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U122 ( .A0_t (wk[57]), .B0_t (DataIn[57]), .Z0_t (Midori_add_Result_Start[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U121 ( .A0_t (wk[56]), .B0_t (DataIn[56]), .Z0_t (Midori_add_Result_Start[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U120 ( .A0_t (wk[55]), .B0_t (DataIn[55]), .Z0_t (Midori_add_Result_Start[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U119 ( .A0_t (wk[54]), .B0_t (DataIn[54]), .Z0_t (Midori_add_Result_Start[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U118 ( .A0_t (wk[53]), .B0_t (DataIn[53]), .Z0_t (Midori_add_Result_Start[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U117 ( .A0_t (wk[52]), .B0_t (DataIn[52]), .Z0_t (Midori_add_Result_Start[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U116 ( .A0_t (wk[51]), .B0_t (DataIn[51]), .Z0_t (Midori_add_Result_Start[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U115 ( .A0_t (wk[50]), .B0_t (DataIn[50]), .Z0_t (Midori_add_Result_Start[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U114 ( .A0_t (wk[49]), .B0_t (DataIn[49]), .Z0_t (Midori_add_Result_Start[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U113 ( .A0_t (wk[48]), .B0_t (DataIn[48]), .Z0_t (Midori_add_Result_Start[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U112 ( .A0_t (wk[47]), .B0_t (DataIn[47]), .Z0_t (Midori_add_Result_Start[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U111 ( .A0_t (wk[46]), .B0_t (DataIn[46]), .Z0_t (Midori_add_Result_Start[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U110 ( .A0_t (wk[45]), .B0_t (DataIn[45]), .Z0_t (Midori_add_Result_Start[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U109 ( .A0_t (wk[44]), .B0_t (DataIn[44]), .Z0_t (Midori_add_Result_Start[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U108 ( .A0_t (wk[43]), .B0_t (DataIn[43]), .Z0_t (Midori_add_Result_Start[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U107 ( .A0_t (wk[42]), .B0_t (DataIn[42]), .Z0_t (Midori_add_Result_Start[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U106 ( .A0_t (wk[41]), .B0_t (DataIn[41]), .Z0_t (Midori_add_Result_Start[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U105 ( .A0_t (wk[40]), .B0_t (DataIn[40]), .Z0_t (Midori_add_Result_Start[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U104 ( .A0_t (wk[39]), .B0_t (DataIn[39]), .Z0_t (Midori_add_Result_Start[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U103 ( .A0_t (wk[38]), .B0_t (DataIn[38]), .Z0_t (Midori_add_Result_Start[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U102 ( .A0_t (wk[37]), .B0_t (DataIn[37]), .Z0_t (Midori_add_Result_Start[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U101 ( .A0_t (wk[36]), .B0_t (DataIn[36]), .Z0_t (Midori_add_Result_Start[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U100 ( .A0_t (wk[35]), .B0_t (DataIn[35]), .Z0_t (Midori_add_Result_Start[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U99 ( .A0_t (wk[34]), .B0_t (DataIn[34]), .Z0_t (Midori_add_Result_Start[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U98 ( .A0_t (wk[33]), .B0_t (DataIn[33]), .Z0_t (Midori_add_Result_Start[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U97 ( .A0_t (wk[32]), .B0_t (DataIn[32]), .Z0_t (Midori_add_Result_Start[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U96 ( .A0_t (wk[31]), .B0_t (DataIn[31]), .Z0_t (Midori_add_Result_Start[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U95 ( .A0_t (wk[30]), .B0_t (DataIn[30]), .Z0_t (Midori_add_Result_Start[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U94 ( .A0_t (wk[29]), .B0_t (DataIn[29]), .Z0_t (Midori_add_Result_Start[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U93 ( .A0_t (wk[28]), .B0_t (DataIn[28]), .Z0_t (Midori_add_Result_Start[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U92 ( .A0_t (wk[27]), .B0_t (DataIn[27]), .Z0_t (Midori_add_Result_Start[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U91 ( .A0_t (wk[26]), .B0_t (DataIn[26]), .Z0_t (Midori_add_Result_Start[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U90 ( .A0_t (wk[25]), .B0_t (DataIn[25]), .Z0_t (Midori_add_Result_Start[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U89 ( .A0_t (wk[24]), .B0_t (DataIn[24]), .Z0_t (Midori_add_Result_Start[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U88 ( .A0_t (wk[23]), .B0_t (DataIn[23]), .Z0_t (Midori_add_Result_Start[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U87 ( .A0_t (wk[22]), .B0_t (DataIn[22]), .Z0_t (Midori_add_Result_Start[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U86 ( .A0_t (wk[21]), .B0_t (DataIn[21]), .Z0_t (Midori_add_Result_Start[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U85 ( .A0_t (wk[20]), .B0_t (DataIn[20]), .Z0_t (Midori_add_Result_Start[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U84 ( .A0_t (wk[19]), .B0_t (DataIn[19]), .Z0_t (Midori_add_Result_Start[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U83 ( .A0_t (wk[18]), .B0_t (DataIn[18]), .Z0_t (Midori_add_Result_Start[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U82 ( .A0_t (wk[17]), .B0_t (DataIn[17]), .Z0_t (Midori_add_Result_Start[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U81 ( .A0_t (wk[16]), .B0_t (DataIn[16]), .Z0_t (Midori_add_Result_Start[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U80 ( .A0_t (wk[15]), .B0_t (DataIn[15]), .Z0_t (Midori_add_Result_Start[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U79 ( .A0_t (wk[14]), .B0_t (DataIn[14]), .Z0_t (Midori_add_Result_Start[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U78 ( .A0_t (wk[13]), .B0_t (DataIn[13]), .Z0_t (Midori_add_Result_Start[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U77 ( .A0_t (wk[12]), .B0_t (DataIn[12]), .Z0_t (Midori_add_Result_Start[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U76 ( .A0_t (wk[11]), .B0_t (DataIn[11]), .Z0_t (Midori_add_Result_Start[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U75 ( .A0_t (wk[10]), .B0_t (DataIn[10]), .Z0_t (Midori_add_Result_Start[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U74 ( .A0_t (wk[9]), .B0_t (DataIn[9]), .Z0_t (Midori_add_Result_Start[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U73 ( .A0_t (wk[8]), .B0_t (DataIn[8]), .Z0_t (Midori_add_Result_Start[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U72 ( .A0_t (wk[7]), .B0_t (DataIn[7]), .Z0_t (Midori_add_Result_Start[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U71 ( .A0_t (wk[6]), .B0_t (DataIn[6]), .Z0_t (Midori_add_Result_Start[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U70 ( .A0_t (wk[5]), .B0_t (DataIn[5]), .Z0_t (Midori_add_Result_Start[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U69 ( .A0_t (wk[4]), .B0_t (DataIn[4]), .Z0_t (Midori_add_Result_Start[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U68 ( .A0_t (wk[3]), .B0_t (DataIn[3]), .Z0_t (Midori_add_Result_Start[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U67 ( .A0_t (wk[2]), .B0_t (DataIn[2]), .Z0_t (Midori_add_Result_Start[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U66 ( .A0_t (wk[1]), .B0_t (DataIn[1]), .Z0_t (Midori_add_Result_Start[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U65 ( .A0_t (wk[0]), .B0_t (DataIn[0]), .Z0_t (Midori_add_Result_Start[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U64 ( .A0_t (wk[56]), .B0_t (Midori_rounds_SR_Result[32]), .Z0_t (DataOut[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U63 ( .A0_t (wk[52]), .B0_t (Midori_rounds_SR_Result[4]), .Z0_t (DataOut[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U62 ( .A0_t (wk[36]), .B0_t (Midori_rounds_SR_Result[16]), .Z0_t (DataOut[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U61 ( .A0_t (wk[32]), .B0_t (Midori_rounds_SR_Result[12]), .Z0_t (DataOut[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U60 ( .A0_t (wk[28]), .B0_t (Midori_rounds_SR_Result[0]), .Z0_t (DataOut[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U59 ( .A0_t (wk[0]), .B0_t (Midori_rounds_SR_Result[48]), .Z0_t (DataOut[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U58 ( .A0_t (wk[59]), .B0_t (Midori_rounds_SR_Result[35]), .Z0_t (DataOut[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U57 ( .A0_t (wk[55]), .B0_t (Midori_rounds_SR_Result[7]), .Z0_t (DataOut[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U56 ( .A0_t (wk[39]), .B0_t (Midori_rounds_SR_Result[19]), .Z0_t (DataOut[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U55 ( .A0_t (wk[35]), .B0_t (Midori_rounds_SR_Result[15]), .Z0_t (DataOut[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U54 ( .A0_t (wk[31]), .B0_t (Midori_rounds_SR_Result[3]), .Z0_t (DataOut[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U53 ( .A0_t (wk[3]), .B0_t (Midori_rounds_SR_Result[51]), .Z0_t (DataOut[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U52 ( .A0_t (wk[63]), .B0_t (Midori_rounds_SR_Result[63]), .Z0_t (DataOut[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U51 ( .A0_t (wk[62]), .B0_t (Midori_rounds_SR_Result[62]), .Z0_t (DataOut[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U50 ( .A0_t (wk[61]), .B0_t (Midori_rounds_SR_Result[61]), .Z0_t (DataOut[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U49 ( .A0_t (wk[58]), .B0_t (Midori_rounds_SR_Result[34]), .Z0_t (DataOut[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U48 ( .A0_t (wk[57]), .B0_t (Midori_rounds_SR_Result[33]), .Z0_t (DataOut[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U47 ( .A0_t (wk[54]), .B0_t (Midori_rounds_SR_Result[6]), .Z0_t (DataOut[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U46 ( .A0_t (wk[53]), .B0_t (Midori_rounds_SR_Result[5]), .Z0_t (DataOut[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U45 ( .A0_t (wk[51]), .B0_t (Midori_rounds_SR_Result[27]), .Z0_t (DataOut[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U44 ( .A0_t (wk[50]), .B0_t (Midori_rounds_SR_Result[26]), .Z0_t (DataOut[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U43 ( .A0_t (wk[49]), .B0_t (Midori_rounds_SR_Result[25]), .Z0_t (DataOut[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U42 ( .A0_t (wk[47]), .B0_t (Midori_rounds_SR_Result[43]), .Z0_t (DataOut[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U41 ( .A0_t (wk[46]), .B0_t (Midori_rounds_SR_Result[42]), .Z0_t (DataOut[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U40 ( .A0_t (wk[45]), .B0_t (Midori_rounds_SR_Result[41]), .Z0_t (DataOut[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U39 ( .A0_t (wk[43]), .B0_t (Midori_rounds_SR_Result[55]), .Z0_t (DataOut[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U38 ( .A0_t (wk[41]), .B0_t (Midori_rounds_SR_Result[53]), .Z0_t (DataOut[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U37 ( .A0_t (wk[38]), .B0_t (Midori_rounds_SR_Result[18]), .Z0_t (DataOut[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U36 ( .A0_t (wk[6]), .B0_t (Midori_rounds_SR_Result[46]), .Z0_t (DataOut[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U35 ( .A0_t (wk[5]), .B0_t (Midori_rounds_SR_Result[45]), .Z0_t (DataOut[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U34 ( .A0_t (wk[2]), .B0_t (Midori_rounds_SR_Result[50]), .Z0_t (DataOut[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U33 ( .A0_t (wk[1]), .B0_t (Midori_rounds_SR_Result[49]), .Z0_t (DataOut[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U32 ( .A0_t (wk[60]), .B0_t (Midori_rounds_SR_Result[60]), .Z0_t (DataOut[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U31 ( .A0_t (wk[48]), .B0_t (Midori_rounds_SR_Result[24]), .Z0_t (DataOut[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U30 ( .A0_t (wk[44]), .B0_t (Midori_rounds_SR_Result[40]), .Z0_t (DataOut[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U29 ( .A0_t (wk[42]), .B0_t (Midori_rounds_SR_Result[54]), .Z0_t (DataOut[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U28 ( .A0_t (wk[37]), .B0_t (Midori_rounds_SR_Result[17]), .Z0_t (DataOut[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U27 ( .A0_t (wk[34]), .B0_t (Midori_rounds_SR_Result[14]), .Z0_t (DataOut[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U26 ( .A0_t (wk[33]), .B0_t (Midori_rounds_SR_Result[13]), .Z0_t (DataOut[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U25 ( .A0_t (wk[30]), .B0_t (Midori_rounds_SR_Result[2]), .Z0_t (DataOut[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U24 ( .A0_t (wk[29]), .B0_t (Midori_rounds_SR_Result[1]), .Z0_t (DataOut[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U23 ( .A0_t (wk[27]), .B0_t (Midori_rounds_SR_Result[31]), .Z0_t (DataOut[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U22 ( .A0_t (wk[26]), .B0_t (Midori_rounds_SR_Result[30]), .Z0_t (DataOut[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U21 ( .A0_t (wk[25]), .B0_t (Midori_rounds_SR_Result[29]), .Z0_t (DataOut[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U20 ( .A0_t (wk[23]), .B0_t (Midori_rounds_SR_Result[59]), .Z0_t (DataOut[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U19 ( .A0_t (wk[22]), .B0_t (Midori_rounds_SR_Result[58]), .Z0_t (DataOut[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U18 ( .A0_t (wk[21]), .B0_t (Midori_rounds_SR_Result[57]), .Z0_t (DataOut[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U17 ( .A0_t (wk[19]), .B0_t (Midori_rounds_SR_Result[39]), .Z0_t (DataOut[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U16 ( .A0_t (wk[18]), .B0_t (Midori_rounds_SR_Result[38]), .Z0_t (DataOut[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U15 ( .A0_t (wk[17]), .B0_t (Midori_rounds_SR_Result[37]), .Z0_t (DataOut[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U14 ( .A0_t (wk[15]), .B0_t (Midori_rounds_SR_Result[23]), .Z0_t (DataOut[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U13 ( .A0_t (wk[14]), .B0_t (Midori_rounds_SR_Result[22]), .Z0_t (DataOut[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U12 ( .A0_t (wk[13]), .B0_t (Midori_rounds_SR_Result[21]), .Z0_t (DataOut[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U11 ( .A0_t (wk[11]), .B0_t (Midori_rounds_SR_Result[11]), .Z0_t (DataOut[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U10 ( .A0_t (wk[10]), .B0_t (Midori_rounds_SR_Result[10]), .Z0_t (DataOut[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U9 ( .A0_t (wk[9]), .B0_t (Midori_rounds_SR_Result[9]), .Z0_t (DataOut[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U8 ( .A0_t (wk[7]), .B0_t (Midori_rounds_SR_Result[47]), .Z0_t (DataOut[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U7 ( .A0_t (wk[40]), .B0_t (Midori_rounds_SR_Result[52]), .Z0_t (DataOut[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U6 ( .A0_t (wk[24]), .B0_t (Midori_rounds_SR_Result[28]), .Z0_t (DataOut[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U5 ( .A0_t (wk[20]), .B0_t (Midori_rounds_SR_Result[56]), .Z0_t (DataOut[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U4 ( .A0_t (wk[16]), .B0_t (Midori_rounds_SR_Result[36]), .Z0_t (DataOut[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U3 ( .A0_t (wk[12]), .B0_t (Midori_rounds_SR_Result[20]), .Z0_t (DataOut[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U2 ( .A0_t (wk[8]), .B0_t (Midori_rounds_SR_Result[8]), .Z0_t (DataOut[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_U1 ( .A0_t (wk[4]), .B0_t (Midori_rounds_SR_Result[44]), .Z0_t (DataOut[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U144 ( .A0_t (Midori_rounds_SR_Result[60]), .B0_t (Midori_rounds_n16), .Z0_t (Midori_rounds_sub_ResultXORkey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U143 ( .A0_t (Midori_rounds_SR_Inv_Result[60]), .B0_t (Midori_rounds_n16), .Z0_t (Midori_rounds_mul_ResultXORkey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U142 ( .A0_t (Midori_rounds_round_Constant[15]), .B0_t (Midori_rounds_SelectedKey[60]), .Z0_t (Midori_rounds_n16) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U141 ( .A0_t (Midori_rounds_SR_Result[44]), .B0_t (Midori_rounds_n15), .Z0_t (Midori_rounds_sub_ResultXORkey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U140 ( .A0_t (Midori_rounds_SR_Inv_Result[52]), .B0_t (Midori_rounds_n15), .Z0_t (Midori_rounds_mul_ResultXORkey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U139 ( .A0_t (Midori_rounds_round_Constant[1]), .B0_t (Midori_rounds_SelectedKey[4]), .Z0_t (Midori_rounds_n15) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U138 ( .A0_t (Midori_rounds_SR_Result[32]), .B0_t (Midori_rounds_n14), .Z0_t (Midori_rounds_sub_ResultXORkey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U137 ( .A0_t (Midori_rounds_SR_Inv_Result[20]), .B0_t (Midori_rounds_n14), .Z0_t (Midori_rounds_mul_ResultXORkey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U136 ( .A0_t (Midori_rounds_round_Constant[14]), .B0_t (Midori_rounds_SelectedKey[56]), .Z0_t (Midori_rounds_n14) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U135 ( .A0_t (Midori_rounds_SR_Result[4]), .B0_t (Midori_rounds_n13), .Z0_t (Midori_rounds_sub_ResultXORkey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U134 ( .A0_t (Midori_rounds_SR_Inv_Result[40]), .B0_t (Midori_rounds_n13), .Z0_t (Midori_rounds_mul_ResultXORkey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U133 ( .A0_t (Midori_rounds_round_Constant[13]), .B0_t (Midori_rounds_SelectedKey[52]), .Z0_t (Midori_rounds_n13) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U132 ( .A0_t (Midori_rounds_SR_Result[20]), .B0_t (Midori_rounds_n12), .Z0_t (Midori_rounds_sub_ResultXORkey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U131 ( .A0_t (Midori_rounds_SR_Inv_Result[32]), .B0_t (Midori_rounds_n12), .Z0_t (Midori_rounds_mul_ResultXORkey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U130 ( .A0_t (Midori_rounds_round_Constant[3]), .B0_t (Midori_rounds_SelectedKey[12]), .Z0_t (Midori_rounds_n12) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U129 ( .A0_t (Midori_rounds_SR_Result[16]), .B0_t (Midori_rounds_n11), .Z0_t (Midori_rounds_sub_ResultXORkey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U128 ( .A0_t (Midori_rounds_SR_Inv_Result[16]), .B0_t (Midori_rounds_n11), .Z0_t (Midori_rounds_mul_ResultXORkey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U127 ( .A0_t (Midori_rounds_round_Constant[9]), .B0_t (Midori_rounds_SelectedKey[36]), .Z0_t (Midori_rounds_n11) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U126 ( .A0_t (Midori_rounds_SR_Result[24]), .B0_t (Midori_rounds_n10), .Z0_t (Midori_rounds_sub_ResultXORkey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U125 ( .A0_t (Midori_rounds_SR_Inv_Result[0]), .B0_t (Midori_rounds_n10), .Z0_t (Midori_rounds_mul_ResultXORkey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U124 ( .A0_t (Midori_rounds_round_Constant[12]), .B0_t (Midori_rounds_SelectedKey[48]), .Z0_t (Midori_rounds_n10) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U123 ( .A0_t (Midori_rounds_SR_Result[12]), .B0_t (Midori_rounds_n9), .Z0_t (Midori_rounds_sub_ResultXORkey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U122 ( .A0_t (Midori_rounds_SR_Inv_Result[56]), .B0_t (Midori_rounds_n9), .Z0_t (Midori_rounds_mul_ResultXORkey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U121 ( .A0_t (Midori_rounds_round_Constant[8]), .B0_t (Midori_rounds_SelectedKey[32]), .Z0_t (Midori_rounds_n9) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U120 ( .A0_t (Midori_rounds_SR_Result[0]), .B0_t (Midori_rounds_n8), .Z0_t (Midori_rounds_sub_ResultXORkey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U119 ( .A0_t (Midori_rounds_SR_Inv_Result[24]), .B0_t (Midori_rounds_n8), .Z0_t (Midori_rounds_mul_ResultXORkey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U118 ( .A0_t (Midori_rounds_round_Constant[7]), .B0_t (Midori_rounds_SelectedKey[28]), .Z0_t (Midori_rounds_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U117 ( .A0_t (Midori_rounds_SR_Result[40]), .B0_t (Midori_rounds_n7), .Z0_t (Midori_rounds_sub_ResultXORkey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U116 ( .A0_t (Midori_rounds_SR_Inv_Result[4]), .B0_t (Midori_rounds_n7), .Z0_t (Midori_rounds_mul_ResultXORkey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U115 ( .A0_t (Midori_rounds_round_Constant[11]), .B0_t (Midori_rounds_SelectedKey[44]), .Z0_t (Midori_rounds_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U114 ( .A0_t (Midori_rounds_SR_Result[28]), .B0_t (Midori_rounds_n6), .Z0_t (Midori_rounds_sub_ResultXORkey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U113 ( .A0_t (Midori_rounds_SR_Inv_Result[48]), .B0_t (Midori_rounds_n6), .Z0_t (Midori_rounds_mul_ResultXORkey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U112 ( .A0_t (Midori_rounds_round_Constant[6]), .B0_t (Midori_rounds_SelectedKey[24]), .Z0_t (Midori_rounds_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U111 ( .A0_t (Midori_rounds_SR_Result[8]), .B0_t (Midori_rounds_n5), .Z0_t (Midori_rounds_sub_ResultXORkey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U110 ( .A0_t (Midori_rounds_SR_Inv_Result[8]), .B0_t (Midori_rounds_n5), .Z0_t (Midori_rounds_mul_ResultXORkey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U109 ( .A0_t (Midori_rounds_round_Constant[2]), .B0_t (Midori_rounds_SelectedKey[8]), .Z0_t (Midori_rounds_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U108 ( .A0_t (Midori_rounds_SR_Result[48]), .B0_t (Midori_rounds_n4), .Z0_t (Midori_rounds_sub_ResultXORkey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U107 ( .A0_t (Midori_rounds_SR_Inv_Result[28]), .B0_t (Midori_rounds_n4), .Z0_t (Midori_rounds_mul_ResultXORkey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U106 ( .A0_t (Midori_rounds_round_Constant[0]), .B0_t (Midori_rounds_SelectedKey[0]), .Z0_t (Midori_rounds_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U105 ( .A0_t (Midori_rounds_SR_Result[52]), .B0_t (Midori_rounds_n3), .Z0_t (Midori_rounds_sub_ResultXORkey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U104 ( .A0_t (Midori_rounds_SR_Inv_Result[44]), .B0_t (Midori_rounds_n3), .Z0_t (Midori_rounds_mul_ResultXORkey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U103 ( .A0_t (Midori_rounds_round_Constant[10]), .B0_t (Midori_rounds_SelectedKey[40]), .Z0_t (Midori_rounds_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U102 ( .A0_t (Midori_rounds_SR_Result[56]), .B0_t (Midori_rounds_n2), .Z0_t (Midori_rounds_sub_ResultXORkey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U101 ( .A0_t (Midori_rounds_SR_Inv_Result[12]), .B0_t (Midori_rounds_n2), .Z0_t (Midori_rounds_mul_ResultXORkey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U100 ( .A0_t (Midori_rounds_round_Constant[5]), .B0_t (Midori_rounds_SelectedKey[20]), .Z0_t (Midori_rounds_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U99 ( .A0_t (Midori_rounds_SR_Result[36]), .B0_t (Midori_rounds_n1), .Z0_t (Midori_rounds_sub_ResultXORkey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U98 ( .A0_t (Midori_rounds_SR_Inv_Result[36]), .B0_t (Midori_rounds_n1), .Z0_t (Midori_rounds_mul_ResultXORkey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_U97 ( .A0_t (Midori_rounds_round_Constant[4]), .B0_t (Midori_rounds_SelectedKey[16]), .Z0_t (Midori_rounds_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U96 ( .A0_t (Midori_rounds_SelectedKey[51]), .B0_t (Midori_rounds_SR_Result[27]), .Z0_t (Midori_rounds_sub_ResultXORkey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U95 ( .A0_t (Midori_rounds_SelectedKey[54]), .B0_t (Midori_rounds_SR_Result[6]), .Z0_t (Midori_rounds_sub_ResultXORkey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U94 ( .A0_t (Midori_rounds_SelectedKey[49]), .B0_t (Midori_rounds_SR_Result[25]), .Z0_t (Midori_rounds_sub_ResultXORkey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U93 ( .A0_t (Midori_rounds_SelectedKey[39]), .B0_t (Midori_rounds_SR_Result[19]), .Z0_t (Midori_rounds_sub_ResultXORkey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U92 ( .A0_t (Midori_rounds_SelectedKey[37]), .B0_t (Midori_rounds_SR_Result[17]), .Z0_t (Midori_rounds_sub_ResultXORkey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U91 ( .A0_t (Midori_rounds_SelectedKey[19]), .B0_t (Midori_rounds_SR_Result[39]), .Z0_t (Midori_rounds_sub_ResultXORkey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U90 ( .A0_t (Midori_rounds_SelectedKey[17]), .B0_t (Midori_rounds_SR_Result[37]), .Z0_t (Midori_rounds_sub_ResultXORkey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U89 ( .A0_t (Midori_rounds_SelectedKey[34]), .B0_t (Midori_rounds_SR_Result[14]), .Z0_t (Midori_rounds_sub_ResultXORkey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U88 ( .A0_t (Midori_rounds_SelectedKey[18]), .B0_t (Midori_rounds_SR_Result[38]), .Z0_t (Midori_rounds_sub_ResultXORkey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U87 ( .A0_t (Midori_rounds_SelectedKey[55]), .B0_t (Midori_rounds_SR_Result[7]), .Z0_t (Midori_rounds_sub_ResultXORkey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U86 ( .A0_t (Midori_rounds_SelectedKey[50]), .B0_t (Midori_rounds_SR_Result[26]), .Z0_t (Midori_rounds_sub_ResultXORkey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U85 ( .A0_t (Midori_rounds_SelectedKey[53]), .B0_t (Midori_rounds_SR_Result[5]), .Z0_t (Midori_rounds_sub_ResultXORkey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U84 ( .A0_t (Midori_rounds_SelectedKey[35]), .B0_t (Midori_rounds_SR_Result[15]), .Z0_t (Midori_rounds_sub_ResultXORkey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U83 ( .A0_t (Midori_rounds_SelectedKey[38]), .B0_t (Midori_rounds_SR_Result[18]), .Z0_t (Midori_rounds_sub_ResultXORkey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U82 ( .A0_t (Midori_rounds_SelectedKey[33]), .B0_t (Midori_rounds_SR_Result[13]), .Z0_t (Midori_rounds_sub_ResultXORkey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U81 ( .A0_t (Midori_rounds_SelectedKey[23]), .B0_t (Midori_rounds_SR_Result[59]), .Z0_t (Midori_rounds_sub_ResultXORkey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U80 ( .A0_t (Midori_rounds_SelectedKey[22]), .B0_t (Midori_rounds_SR_Result[58]), .Z0_t (Midori_rounds_sub_ResultXORkey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U79 ( .A0_t (Midori_rounds_SelectedKey[21]), .B0_t (Midori_rounds_SR_Result[57]), .Z0_t (Midori_rounds_sub_ResultXORkey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U78 ( .A0_t (Midori_rounds_SelectedKey[7]), .B0_t (Midori_rounds_SR_Result[47]), .Z0_t (Midori_rounds_sub_ResultXORkey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U77 ( .A0_t (Midori_rounds_SelectedKey[2]), .B0_t (Midori_rounds_SR_Result[50]), .Z0_t (Midori_rounds_sub_ResultXORkey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U76 ( .A0_t (Midori_rounds_SelectedKey[5]), .B0_t (Midori_rounds_SR_Result[45]), .Z0_t (Midori_rounds_sub_ResultXORkey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U75 ( .A0_t (Midori_rounds_SelectedKey[3]), .B0_t (Midori_rounds_SR_Result[51]), .Z0_t (Midori_rounds_sub_ResultXORkey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U74 ( .A0_t (Midori_rounds_SelectedKey[6]), .B0_t (Midori_rounds_SR_Result[46]), .Z0_t (Midori_rounds_sub_ResultXORkey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U73 ( .A0_t (Midori_rounds_SelectedKey[1]), .B0_t (Midori_rounds_SR_Result[49]), .Z0_t (Midori_rounds_sub_ResultXORkey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U72 ( .A0_t (Midori_rounds_SelectedKey[63]), .B0_t (Midori_rounds_SR_Inv_Result[63]), .Z0_t (Midori_rounds_mul_ResultXORkey[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U71 ( .A0_t (Midori_rounds_SelectedKey[62]), .B0_t (Midori_rounds_SR_Inv_Result[62]), .Z0_t (Midori_rounds_mul_ResultXORkey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U70 ( .A0_t (Midori_rounds_SelectedKey[61]), .B0_t (Midori_rounds_SR_Inv_Result[61]), .Z0_t (Midori_rounds_mul_ResultXORkey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U69 ( .A0_t (Midori_rounds_SelectedKey[59]), .B0_t (Midori_rounds_SR_Inv_Result[23]), .Z0_t (Midori_rounds_mul_ResultXORkey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U68 ( .A0_t (Midori_rounds_SelectedKey[58]), .B0_t (Midori_rounds_SR_Inv_Result[22]), .Z0_t (Midori_rounds_mul_ResultXORkey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U67 ( .A0_t (Midori_rounds_SelectedKey[57]), .B0_t (Midori_rounds_SR_Inv_Result[21]), .Z0_t (Midori_rounds_mul_ResultXORkey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U66 ( .A0_t (Midori_rounds_SelectedKey[55]), .B0_t (Midori_rounds_SR_Inv_Result[43]), .Z0_t (Midori_rounds_mul_ResultXORkey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U65 ( .A0_t (Midori_rounds_SelectedKey[54]), .B0_t (Midori_rounds_SR_Inv_Result[42]), .Z0_t (Midori_rounds_mul_ResultXORkey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U64 ( .A0_t (Midori_rounds_SelectedKey[53]), .B0_t (Midori_rounds_SR_Inv_Result[41]), .Z0_t (Midori_rounds_mul_ResultXORkey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U63 ( .A0_t (Midori_rounds_SelectedKey[51]), .B0_t (Midori_rounds_SR_Inv_Result[3]), .Z0_t (Midori_rounds_mul_ResultXORkey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U62 ( .A0_t (Midori_rounds_SelectedKey[50]), .B0_t (Midori_rounds_SR_Inv_Result[2]), .Z0_t (Midori_rounds_mul_ResultXORkey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U61 ( .A0_t (Midori_rounds_SelectedKey[49]), .B0_t (Midori_rounds_SR_Inv_Result[1]), .Z0_t (Midori_rounds_mul_ResultXORkey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U60 ( .A0_t (Midori_rounds_SelectedKey[47]), .B0_t (Midori_rounds_SR_Inv_Result[7]), .Z0_t (Midori_rounds_mul_ResultXORkey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U59 ( .A0_t (Midori_rounds_SelectedKey[46]), .B0_t (Midori_rounds_SR_Inv_Result[6]), .Z0_t (Midori_rounds_mul_ResultXORkey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U58 ( .A0_t (Midori_rounds_SelectedKey[45]), .B0_t (Midori_rounds_SR_Inv_Result[5]), .Z0_t (Midori_rounds_mul_ResultXORkey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U57 ( .A0_t (Midori_rounds_SelectedKey[43]), .B0_t (Midori_rounds_SR_Inv_Result[47]), .Z0_t (Midori_rounds_mul_ResultXORkey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U56 ( .A0_t (Midori_rounds_SelectedKey[42]), .B0_t (Midori_rounds_SR_Inv_Result[46]), .Z0_t (Midori_rounds_mul_ResultXORkey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U55 ( .A0_t (Midori_rounds_SelectedKey[41]), .B0_t (Midori_rounds_SR_Inv_Result[45]), .Z0_t (Midori_rounds_mul_ResultXORkey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U54 ( .A0_t (Midori_rounds_SelectedKey[39]), .B0_t (Midori_rounds_SR_Inv_Result[19]), .Z0_t (Midori_rounds_mul_ResultXORkey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U53 ( .A0_t (Midori_rounds_SelectedKey[38]), .B0_t (Midori_rounds_SR_Inv_Result[18]), .Z0_t (Midori_rounds_mul_ResultXORkey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U52 ( .A0_t (Midori_rounds_SelectedKey[37]), .B0_t (Midori_rounds_SR_Inv_Result[17]), .Z0_t (Midori_rounds_mul_ResultXORkey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U51 ( .A0_t (Midori_rounds_SelectedKey[35]), .B0_t (Midori_rounds_SR_Inv_Result[59]), .Z0_t (Midori_rounds_mul_ResultXORkey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U50 ( .A0_t (Midori_rounds_SelectedKey[34]), .B0_t (Midori_rounds_SR_Inv_Result[58]), .Z0_t (Midori_rounds_mul_ResultXORkey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U49 ( .A0_t (Midori_rounds_SelectedKey[33]), .B0_t (Midori_rounds_SR_Inv_Result[57]), .Z0_t (Midori_rounds_mul_ResultXORkey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U48 ( .A0_t (Midori_rounds_SelectedKey[31]), .B0_t (Midori_rounds_SR_Inv_Result[27]), .Z0_t (Midori_rounds_mul_ResultXORkey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U47 ( .A0_t (Midori_rounds_SelectedKey[30]), .B0_t (Midori_rounds_SR_Inv_Result[26]), .Z0_t (Midori_rounds_mul_ResultXORkey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U46 ( .A0_t (Midori_rounds_SelectedKey[29]), .B0_t (Midori_rounds_SR_Inv_Result[25]), .Z0_t (Midori_rounds_mul_ResultXORkey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U45 ( .A0_t (Midori_rounds_SelectedKey[27]), .B0_t (Midori_rounds_SR_Inv_Result[51]), .Z0_t (Midori_rounds_mul_ResultXORkey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U44 ( .A0_t (Midori_rounds_SelectedKey[26]), .B0_t (Midori_rounds_SR_Inv_Result[50]), .Z0_t (Midori_rounds_mul_ResultXORkey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U43 ( .A0_t (Midori_rounds_SelectedKey[25]), .B0_t (Midori_rounds_SR_Inv_Result[49]), .Z0_t (Midori_rounds_mul_ResultXORkey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U42 ( .A0_t (Midori_rounds_SelectedKey[23]), .B0_t (Midori_rounds_SR_Inv_Result[15]), .Z0_t (Midori_rounds_mul_ResultXORkey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U41 ( .A0_t (Midori_rounds_SelectedKey[22]), .B0_t (Midori_rounds_SR_Inv_Result[14]), .Z0_t (Midori_rounds_mul_ResultXORkey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U40 ( .A0_t (Midori_rounds_SelectedKey[21]), .B0_t (Midori_rounds_SR_Inv_Result[13]), .Z0_t (Midori_rounds_mul_ResultXORkey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U39 ( .A0_t (Midori_rounds_SelectedKey[19]), .B0_t (Midori_rounds_SR_Inv_Result[39]), .Z0_t (Midori_rounds_mul_ResultXORkey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U38 ( .A0_t (Midori_rounds_SelectedKey[18]), .B0_t (Midori_rounds_SR_Inv_Result[38]), .Z0_t (Midori_rounds_mul_ResultXORkey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U37 ( .A0_t (Midori_rounds_SelectedKey[17]), .B0_t (Midori_rounds_SR_Inv_Result[37]), .Z0_t (Midori_rounds_mul_ResultXORkey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U36 ( .A0_t (Midori_rounds_SelectedKey[15]), .B0_t (Midori_rounds_SR_Inv_Result[35]), .Z0_t (Midori_rounds_mul_ResultXORkey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U35 ( .A0_t (Midori_rounds_SelectedKey[14]), .B0_t (Midori_rounds_SR_Inv_Result[34]), .Z0_t (Midori_rounds_mul_ResultXORkey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U34 ( .A0_t (Midori_rounds_SelectedKey[13]), .B0_t (Midori_rounds_SR_Inv_Result[33]), .Z0_t (Midori_rounds_mul_ResultXORkey[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U33 ( .A0_t (Midori_rounds_SelectedKey[11]), .B0_t (Midori_rounds_SR_Inv_Result[11]), .Z0_t (Midori_rounds_mul_ResultXORkey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U32 ( .A0_t (Midori_rounds_SelectedKey[10]), .B0_t (Midori_rounds_SR_Inv_Result[10]), .Z0_t (Midori_rounds_mul_ResultXORkey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U31 ( .A0_t (Midori_rounds_SelectedKey[9]), .B0_t (Midori_rounds_SR_Inv_Result[9]), .Z0_t (Midori_rounds_mul_ResultXORkey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U30 ( .A0_t (Midori_rounds_SelectedKey[7]), .B0_t (Midori_rounds_SR_Inv_Result[55]), .Z0_t (Midori_rounds_mul_ResultXORkey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U29 ( .A0_t (Midori_rounds_SelectedKey[6]), .B0_t (Midori_rounds_SR_Inv_Result[54]), .Z0_t (Midori_rounds_mul_ResultXORkey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U28 ( .A0_t (Midori_rounds_SelectedKey[5]), .B0_t (Midori_rounds_SR_Inv_Result[53]), .Z0_t (Midori_rounds_mul_ResultXORkey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U27 ( .A0_t (Midori_rounds_SelectedKey[3]), .B0_t (Midori_rounds_SR_Inv_Result[31]), .Z0_t (Midori_rounds_mul_ResultXORkey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U26 ( .A0_t (Midori_rounds_SelectedKey[2]), .B0_t (Midori_rounds_SR_Inv_Result[30]), .Z0_t (Midori_rounds_mul_ResultXORkey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U25 ( .A0_t (Midori_rounds_SelectedKey[1]), .B0_t (Midori_rounds_SR_Inv_Result[29]), .Z0_t (Midori_rounds_mul_ResultXORkey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U24 ( .A0_t (Midori_rounds_SelectedKey[43]), .B0_t (Midori_rounds_SR_Result[55]), .Z0_t (Midori_rounds_sub_ResultXORkey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U23 ( .A0_t (Midori_rounds_SelectedKey[41]), .B0_t (Midori_rounds_SR_Result[53]), .Z0_t (Midori_rounds_sub_ResultXORkey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U22 ( .A0_t (Midori_rounds_SelectedKey[31]), .B0_t (Midori_rounds_SR_Result[3]), .Z0_t (Midori_rounds_sub_ResultXORkey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U21 ( .A0_t (Midori_rounds_SelectedKey[29]), .B0_t (Midori_rounds_SR_Result[1]), .Z0_t (Midori_rounds_sub_ResultXORkey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U20 ( .A0_t (Midori_rounds_SelectedKey[63]), .B0_t (Midori_rounds_SR_Result[63]), .Z0_t (Midori_rounds_sub_ResultXORkey[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U19 ( .A0_t (Midori_rounds_SelectedKey[61]), .B0_t (Midori_rounds_SR_Result[61]), .Z0_t (Midori_rounds_sub_ResultXORkey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U18 ( .A0_t (Midori_rounds_SelectedKey[26]), .B0_t (Midori_rounds_SR_Result[30]), .Z0_t (Midori_rounds_sub_ResultXORkey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U17 ( .A0_t (Midori_rounds_SelectedKey[62]), .B0_t (Midori_rounds_SR_Result[62]), .Z0_t (Midori_rounds_sub_ResultXORkey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U16 ( .A0_t (Midori_rounds_SelectedKey[42]), .B0_t (Midori_rounds_SR_Result[54]), .Z0_t (Midori_rounds_sub_ResultXORkey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U15 ( .A0_t (Midori_rounds_SelectedKey[59]), .B0_t (Midori_rounds_SR_Result[35]), .Z0_t (Midori_rounds_sub_ResultXORkey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U14 ( .A0_t (Midori_rounds_SelectedKey[58]), .B0_t (Midori_rounds_SR_Result[34]), .Z0_t (Midori_rounds_sub_ResultXORkey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U13 ( .A0_t (Midori_rounds_SelectedKey[57]), .B0_t (Midori_rounds_SR_Result[33]), .Z0_t (Midori_rounds_sub_ResultXORkey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U12 ( .A0_t (Midori_rounds_SelectedKey[47]), .B0_t (Midori_rounds_SR_Result[43]), .Z0_t (Midori_rounds_sub_ResultXORkey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U11 ( .A0_t (Midori_rounds_SelectedKey[46]), .B0_t (Midori_rounds_SR_Result[42]), .Z0_t (Midori_rounds_sub_ResultXORkey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U10 ( .A0_t (Midori_rounds_SelectedKey[45]), .B0_t (Midori_rounds_SR_Result[41]), .Z0_t (Midori_rounds_sub_ResultXORkey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U9 ( .A0_t (Midori_rounds_SelectedKey[27]), .B0_t (Midori_rounds_SR_Result[31]), .Z0_t (Midori_rounds_sub_ResultXORkey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U8 ( .A0_t (Midori_rounds_SelectedKey[30]), .B0_t (Midori_rounds_SR_Result[2]), .Z0_t (Midori_rounds_sub_ResultXORkey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U7 ( .A0_t (Midori_rounds_SelectedKey[25]), .B0_t (Midori_rounds_SR_Result[29]), .Z0_t (Midori_rounds_sub_ResultXORkey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U6 ( .A0_t (Midori_rounds_SelectedKey[11]), .B0_t (Midori_rounds_SR_Result[11]), .Z0_t (Midori_rounds_sub_ResultXORkey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U5 ( .A0_t (Midori_rounds_SelectedKey[10]), .B0_t (Midori_rounds_SR_Result[10]), .Z0_t (Midori_rounds_sub_ResultXORkey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U4 ( .A0_t (Midori_rounds_SelectedKey[9]), .B0_t (Midori_rounds_SR_Result[9]), .Z0_t (Midori_rounds_sub_ResultXORkey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U3 ( .A0_t (Midori_rounds_SelectedKey[15]), .B0_t (Midori_rounds_SR_Result[23]), .Z0_t (Midori_rounds_sub_ResultXORkey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U2 ( .A0_t (Midori_rounds_SelectedKey[14]), .B0_t (Midori_rounds_SR_Result[22]), .Z0_t (Midori_rounds_sub_ResultXORkey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_U1 ( .A0_t (Midori_rounds_SelectedKey[13]), .B0_t (Midori_rounds_SR_Result[21]), .Z0_t (Midori_rounds_sub_ResultXORkey[13]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U134 ( .A0_t (Midori_rounds_constant_MUX_n139), .B0_t (Midori_rounds_constant_MUX_n138), .Z0_t (Midori_rounds_round_Constant[3]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U133 ( .A0_t (Midori_rounds_constant_MUX_n137), .B0_t (Midori_rounds_constant_MUX_n136), .Z0_t (Midori_rounds_constant_MUX_n138) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U132 ( .A0_t (Midori_rounds_constant_MUX_n103), .B0_t (Midori_rounds_constant_MUX_n134), .Z0_t (Midori_rounds_round_Constant[9]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U131 ( .A0_t (Midori_rounds_constant_MUX_n133), .B0_t (Midori_rounds_constant_MUX_n132), .Z0_t (Midori_rounds_constant_MUX_n134) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U130 ( .A0_t (Midori_rounds_constant_MUX_n131), .B0_t (Midori_rounds_constant_MUX_n130), .Z0_t (Midori_rounds_constant_MUX_n132) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U129 ( .A0_t (Midori_rounds_constant_MUX_n129), .B0_t (Midori_rounds_constant_MUX_n128), .Z0_t (Midori_rounds_round_Constant[11]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U128 ( .A0_t (Midori_rounds_constant_MUX_n125), .B0_t (Midori_rounds_constant_MUX_n126), .Z0_t (Midori_rounds_constant_MUX_n128) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U126 ( .A0_t (Midori_rounds_constant_MUX_n124), .B0_t (Midori_rounds_constant_MUX_n123), .Z0_t (Midori_rounds_constant_MUX_n129) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U125 ( .A0_t (Midori_rounds_constant_MUX_n122), .B0_t (Midori_rounds_constant_MUX_n120), .Z0_t (Midori_rounds_constant_MUX_n124) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U124 ( .A0_t (Midori_rounds_constant_MUX_n119), .B0_t (Midori_rounds_constant_MUX_n118), .Z0_t (Midori_rounds_constant_MUX_n122) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U123 ( .A0_t (Midori_rounds_constant_MUX_n117), .B0_t (Midori_rounds_constant_MUX_n116), .Z0_t (Midori_rounds_round_Constant[12]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U122 ( .A0_t (Midori_rounds_constant_MUX_n115), .B0_t (Midori_rounds_constant_MUX_n114), .Z0_t (Midori_rounds_constant_MUX_n116) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U121 ( .A0_t (Midori_rounds_constant_MUX_n113), .B0_t (Midori_rounds_constant_MUX_n110), .Z0_t (Midori_rounds_round_Constant[7]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U120 ( .A0_t (Midori_rounds_constant_MUX_n109), .B0_t (Midori_rounds_constant_MUX_n108), .Z0_t (Midori_rounds_constant_MUX_n110) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U118 ( .A0_t (Midori_rounds_constant_MUX_n133), .B0_t (Midori_rounds_constant_MUX_n115), .Z0_t (Midori_rounds_constant_MUX_n113) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U117 ( .A0_t (Midori_rounds_constant_MUX_n103), .B0_t (Midori_rounds_constant_MUX_n107), .Z0_t (Midori_rounds_round_Constant[15]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U116 ( .A0_t (Midori_rounds_constant_MUX_n136), .B0_t (Midori_rounds_constant_MUX_n106), .Z0_t (Midori_rounds_constant_MUX_n107) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U115 ( .A0_t (Midori_rounds_constant_MUX_n83), .B0_t (Midori_rounds_constant_MUX_n104), .Z0_t (Midori_rounds_constant_MUX_n106) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U113 ( .A0_t (Midori_rounds_constant_MUX_n102), .B0_t (Midori_rounds_constant_MUX_n130), .Z0_t (Midori_rounds_round_Constant[14]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U112 ( .A0_t (Midori_rounds_constant_MUX_n101), .B0_t (Midori_rounds_constant_MUX_n108), .Z0_t (Midori_rounds_constant_MUX_n102) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U111 ( .A0_t (Midori_rounds_constant_MUX_n100), .B0_t (Midori_rounds_constant_MUX_n99), .Z0_t (Midori_rounds_constant_MUX_n108) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U110 ( .A0_t (Midori_rounds_constant_MUX_n103), .B0_t (Midori_rounds_constant_MUX_n137), .Z0_t (Midori_rounds_constant_MUX_n99) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U109 ( .A0_t (Midori_rounds_constant_MUX_n98), .B0_t (Midori_rounds_constant_MUX_n97), .Z0_t (Midori_rounds_round_Constant[10]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U108 ( .A0_t (Midori_rounds_constant_MUX_n96), .B0_t (Midori_rounds_constant_MUX_n95), .Z0_t (Midori_rounds_constant_MUX_n98) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U107 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_constant_MUX_n94), .Z0_t (Midori_rounds_constant_MUX_n95) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U106 ( .A0_t (Midori_rounds_constant_MUX_n93), .B0_t (Midori_rounds_constant_MUX_n92), .Z0_t (Midori_rounds_constant_MUX_n94) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U105 ( .A0_t (Midori_rounds_constant_MUX_n118), .B0_t (Midori_rounds_constant_MUX_n91), .Z0_t (Midori_rounds_constant_MUX_n92) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U104 ( .A0_t (enc_dec), .B0_t (Midori_rounds_constant_MUX_n123), .Z0_t (Midori_rounds_constant_MUX_n91) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U103 ( .A0_t (Midori_rounds_constant_MUX_n35), .B0_t (Midori_rounds_constant_MUX_n88), .Z0_t (Midori_rounds_constant_MUX_n123) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U102 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n86), .Z0_t (Midori_rounds_constant_MUX_n118) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U101 ( .A0_t (Midori_rounds_constant_MUX_n85), .B0_t (Midori_rounds_constant_MUX_n125), .Z0_t (Midori_rounds_round_Constant[6]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U100 ( .A0_t (Midori_rounds_constant_MUX_n114), .B0_t (Midori_rounds_constant_MUX_n84), .Z0_t (Midori_rounds_constant_MUX_n85) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U99 ( .A0_t (Midori_rounds_constant_MUX_n83), .B0_t (Midori_rounds_constant_MUX_n131), .Z0_t (Midori_rounds_constant_MUX_n84) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U97 ( .A0_t (Midori_rounds_constant_MUX_n82), .B0_t (Midori_rounds_constant_MUX_n81), .Z0_t (Midori_rounds_constant_MUX_n114) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U96 ( .A0_t (Midori_rounds_constant_MUX_n80), .B0_t (Midori_rounds_constant_MUX_n79), .Z0_t (Midori_rounds_round_Constant[5]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U95 ( .A0_t (Midori_rounds_constant_MUX_n137), .B0_t (Midori_rounds_constant_MUX_n78), .Z0_t (Midori_rounds_constant_MUX_n79) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U94 ( .A0_t (Midori_rounds_constant_MUX_n77), .B0_t (Midori_rounds_constant_MUX_n76), .Z0_t (Midori_rounds_round_Constant[1]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U93 ( .A0_t (Midori_rounds_constant_MUX_n136), .B0_t (Midori_rounds_constant_MUX_n75), .Z0_t (Midori_rounds_constant_MUX_n77) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U92 ( .A0_t (Midori_rounds_constant_MUX_n74), .B0_t (Midori_rounds_constant_MUX_n131), .Z0_t (Midori_rounds_constant_MUX_n75) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U91 ( .A0_t (Midori_rounds_constant_MUX_n73), .B0_t (Midori_rounds_constant_MUX_n72), .Z0_t (Midori_rounds_constant_MUX_n136) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U90 ( .A0_t (Midori_rounds_constant_MUX_n126), .B0_t (enc_dec), .Z0_t (Midori_rounds_constant_MUX_n72) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U88 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_constant_MUX_n70), .Z0_t (Midori_rounds_constant_MUX_n126) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U87 ( .A0_t (Midori_rounds_constant_MUX_n69), .B0_t (Midori_rounds_constant_MUX_n111), .Z0_t (Midori_rounds_constant_MUX_n73) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U86 ( .A0_t (Midori_rounds_constant_MUX_n100), .B0_t (Midori_rounds_constant_MUX_n68), .Z0_t (Midori_rounds_round_Constant[13]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U85 ( .A0_t (Midori_rounds_constant_MUX_n76), .B0_t (Midori_rounds_constant_MUX_n66), .Z0_t (Midori_rounds_constant_MUX_n68) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U83 ( .A0_t (Midori_rounds_constant_MUX_n42), .B0_t (Midori_rounds_constant_MUX_n82), .Z0_t (Midori_rounds_constant_MUX_n100) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U82 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_constant_MUX_n64), .Z0_t (Midori_rounds_constant_MUX_n82) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U81 ( .A0_t (Midori_rounds_constant_MUX_n70), .B0_t (Midori_rounds_constant_MUX_n62), .Z0_t (Midori_rounds_constant_MUX_n64) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U80 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n69), .Z0_t (Midori_rounds_constant_MUX_n62) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U79 ( .A0_t (Midori_rounds_constant_MUX_n117), .B0_t (Midori_rounds_constant_MUX_n61), .Z0_t (Midori_rounds_round_Constant[4]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U78 ( .A0_t (Midori_rounds_constant_MUX_n137), .B0_t (Midori_rounds_constant_MUX_n66), .Z0_t (Midori_rounds_constant_MUX_n61) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U77 ( .A0_t (Midori_rounds_constant_MUX_n60), .B0_t (Midori_rounds_constant_MUX_n130), .Z0_t (Midori_rounds_constant_MUX_n66) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U76 ( .A0_t (Midori_rounds_constant_MUX_n59), .B0_t (Midori_rounds_constant_MUX_n58), .Z0_t (Midori_rounds_constant_MUX_n137) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U75 ( .A0_t (Midori_rounds_constant_MUX_n88), .B0_t (Midori_rounds_constant_MUX_n121), .Z0_t (Midori_rounds_constant_MUX_n58) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U74 ( .A0_t (Midori_rounds_constant_MUX_n57), .B0_t (Midori_rounds_constant_MUX_n56), .Z0_t (Midori_rounds_constant_MUX_n59) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U73 ( .A0_t (Midori_rounds_constant_MUX_n55), .B0_t (round_Signal[2]), .Z0_t (Midori_rounds_constant_MUX_n121) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U72 ( .A0_t (Midori_rounds_constant_MUX_n139), .B0_t (Midori_rounds_constant_MUX_n54), .Z0_t (Midori_rounds_round_Constant[2]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U71 ( .A0_t (Midori_rounds_constant_MUX_n42), .B0_t (Midori_rounds_constant_MUX_n78), .Z0_t (Midori_rounds_constant_MUX_n54) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U70 ( .A0_t (Midori_rounds_constant_MUX_n60), .B0_t (Midori_rounds_constant_MUX_n131), .Z0_t (Midori_rounds_constant_MUX_n78) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U69 ( .A0_t (Midori_rounds_constant_MUX_n53), .B0_t (Midori_rounds_constant_MUX_n52), .Z0_t (Midori_rounds_constant_MUX_n131) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U68 ( .A0_t (Midori_rounds_constant_MUX_n119), .B0_t (Midori_rounds_constant_MUX_n51), .Z0_t (Midori_rounds_constant_MUX_n52) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U67 ( .A0_t (Midori_rounds_constant_MUX_n88), .B0_t (Midori_rounds_constant_MUX_n50), .Z0_t (Midori_rounds_constant_MUX_n53) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U66 ( .A0_t (Midori_rounds_constant_MUX_n133), .B0_t (Midori_rounds_constant_MUX_n81), .Z0_t (Midori_rounds_constant_MUX_n139) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U65 ( .A0_t (Midori_rounds_constant_MUX_n125), .B0_t (Midori_rounds_constant_MUX_n76), .Z0_t (Midori_rounds_constant_MUX_n133) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U64 ( .A0_t (round_Signal[1]), .B0_t (Midori_rounds_constant_MUX_n112), .Z0_t (Midori_rounds_constant_MUX_n76) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U63 ( .A0_t (Midori_rounds_constant_MUX_n104), .B0_t (Midori_rounds_constant_MUX_n74), .Z0_t (Midori_rounds_round_Constant[0]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U62 ( .A0_t (Midori_rounds_constant_MUX_n109), .B0_t (Midori_rounds_constant_MUX_n49), .Z0_t (Midori_rounds_constant_MUX_n74) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U61 ( .A0_t (Midori_rounds_constant_MUX_n48), .B0_t (Midori_rounds_constant_MUX_n130), .Z0_t (Midori_rounds_constant_MUX_n49) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U60 ( .A0_t (round_Signal[1]), .B0_t (Midori_rounds_constant_MUX_n43), .Z0_t (Midori_rounds_constant_MUX_n130) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U59 ( .A0_t (Midori_rounds_constant_MUX_n42), .B0_t (Midori_rounds_constant_MUX_n81), .Z0_t (Midori_rounds_constant_MUX_n48) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U58 ( .A0_t (Midori_rounds_constant_MUX_n47), .B0_t (Midori_rounds_constant_MUX_n46), .Z0_t (Midori_rounds_constant_MUX_n81) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U57 ( .A0_t (Midori_rounds_constant_MUX_n86), .B0_t (Midori_rounds_constant_MUX_n50), .Z0_t (Midori_rounds_constant_MUX_n46) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U55 ( .A0_t (Midori_rounds_constant_MUX_n57), .B0_t (Midori_rounds_constant_MUX_n119), .Z0_t (Midori_rounds_constant_MUX_n47) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U52 ( .A0_t (Midori_rounds_constant_MUX_n60), .B0_t (Midori_rounds_constant_MUX_n115), .Z0_t (Midori_rounds_constant_MUX_n104) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U51 ( .A0_t (Midori_rounds_constant_MUX_n97), .B0_t (Midori_rounds_constant_MUX_n40), .Z0_t (Midori_rounds_constant_MUX_n115) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U50 ( .A0_t (Midori_rounds_constant_MUX_n88), .B0_t (Midori_rounds_constant_MUX_n36), .Z0_t (Midori_rounds_constant_MUX_n40) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U49 ( .A0_t (Midori_rounds_constant_MUX_n51), .B0_t (Midori_rounds_constant_MUX_n34), .Z0_t (Midori_rounds_constant_MUX_n97) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U47 ( .A0_t (Midori_rounds_constant_MUX_n96), .B0_t (Midori_rounds_constant_MUX_n37), .Z0_t (Midori_rounds_constant_MUX_n60) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U46 ( .A0_t (Midori_rounds_constant_MUX_n36), .B0_t (Midori_rounds_constant_MUX_n35), .Z0_t (Midori_rounds_constant_MUX_n37) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U45 ( .A0_t (Midori_rounds_constant_MUX_n34), .B0_t (Midori_rounds_constant_MUX_n70), .Z0_t (Midori_rounds_constant_MUX_n96) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U44 ( .A0_t (Midori_rounds_constant_MUX_n117), .B0_t (Midori_rounds_constant_MUX_n125), .Z0_t (Midori_rounds_round_Constant[8]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U43 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_constant_MUX_n51), .Z0_t (Midori_rounds_constant_MUX_n125) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U42 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n35), .Z0_t (Midori_rounds_constant_MUX_n51) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U41 ( .A0_t (Midori_rounds_constant_MUX_n103), .B0_t (Midori_rounds_constant_MUX_n33), .Z0_t (Midori_rounds_constant_MUX_n117) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U40 ( .A0_t (Midori_rounds_constant_MUX_n80), .B0_t (Midori_rounds_constant_MUX_n42), .Z0_t (Midori_rounds_constant_MUX_n33) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U39 ( .A0_t (Midori_rounds_constant_MUX_n32), .B0_t (Midori_rounds_constant_MUX_n31), .Z0_t (Midori_rounds_constant_MUX_n42) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U38 ( .A0_t (Midori_rounds_constant_MUX_n57), .B0_t (Midori_rounds_constant_MUX_n34), .Z0_t (Midori_rounds_constant_MUX_n31) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U37 ( .A0_t (Midori_rounds_constant_MUX_n86), .B0_t (Midori_rounds_constant_MUX_n36), .Z0_t (Midori_rounds_constant_MUX_n32) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U36 ( .A0_t (Midori_rounds_constant_MUX_n101), .B0_t (Midori_rounds_constant_MUX_n109), .Z0_t (Midori_rounds_constant_MUX_n80) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U35 ( .A0_t (Midori_rounds_constant_MUX_n30), .B0_t (Midori_rounds_constant_MUX_n29), .Z0_t (Midori_rounds_constant_MUX_n109) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U34 ( .A0_t (Midori_rounds_constant_MUX_n93), .B0_t (Midori_rounds_constant_MUX_n34), .Z0_t (Midori_rounds_constant_MUX_n29) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U32 ( .A0_t (Midori_rounds_constant_MUX_n36), .B0_t (Midori_rounds_constant_MUX_n69), .Z0_t (Midori_rounds_constant_MUX_n30) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U30 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n119), .Z0_t (Midori_rounds_constant_MUX_n36) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U29 ( .A0_t (Midori_rounds_constant_MUX_n28), .B0_t (Midori_rounds_constant_MUX_n27), .Z0_t (Midori_rounds_constant_MUX_n101) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U28 ( .A0_t (Midori_rounds_constant_MUX_n35), .B0_t (Midori_rounds_constant_MUX_n50), .Z0_t (Midori_rounds_constant_MUX_n27) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U26 ( .A0_t (round_Signal[3]), .B0_t (round_Signal[1]), .Z0_t (Midori_rounds_constant_MUX_n35) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U25 ( .A0_t (Midori_rounds_constant_MUX_n83), .B0_t (Midori_rounds_constant_MUX_n25), .Z0_t (Midori_rounds_constant_MUX_n28) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U24 ( .A0_t (Midori_rounds_constant_MUX_n119), .B0_t (Midori_rounds_constant_MUX_n70), .Z0_t (Midori_rounds_constant_MUX_n25) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U22 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n88), .Z0_t (Midori_rounds_constant_MUX_n70) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U21 ( .A0_t (Midori_rounds_constant_MUX_n24), .B0_t (Midori_rounds_constant_MUX_n23), .Z0_t (Midori_rounds_constant_MUX_n83) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U20 ( .A0_t (Midori_rounds_constant_MUX_n55), .B0_t (Midori_rounds_constant_MUX_n57), .Z0_t (Midori_rounds_constant_MUX_n23) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U18 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n69), .Z0_t (Midori_rounds_constant_MUX_n57) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U17 ( .A0_t (enc_dec), .B0_t (round_Signal[0]), .Z0_t (Midori_rounds_constant_MUX_n55) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U16 ( .A0_t (Midori_rounds_constant_MUX_n111), .B0_t (Midori_rounds_constant_MUX_n88), .Z0_t (Midori_rounds_constant_MUX_n24) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U15 ( .A0_t (round_Signal[1]), .B0_t (round_Signal[3]), .Z0_t (Midori_rounds_constant_MUX_n88) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U13 ( .A0_t (Midori_rounds_constant_MUX_n22), .B0_t (Midori_rounds_constant_MUX_n120), .Z0_t (Midori_rounds_constant_MUX_n103) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U12 ( .A0_t (Midori_rounds_constant_MUX_n119), .B0_t (Midori_rounds_constant_MUX_n93), .Z0_t (Midori_rounds_constant_MUX_n120) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U11 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n86), .Z0_t (Midori_rounds_constant_MUX_n93) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U10 ( .A0_t (round_Signal[3]), .B0_t (round_Signal[1]), .Z0_t (Midori_rounds_constant_MUX_n86) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U8 ( .A0_t (round_Signal[0]), .B0_t (enc_dec), .Z0_t (Midori_rounds_constant_MUX_n119) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U7 ( .A0_t (Midori_rounds_constant_MUX_n50), .B0_t (Midori_rounds_constant_MUX_n69), .Z0_t (Midori_rounds_constant_MUX_n22) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U6 ( .A0_t (round_Signal[3]), .B0_t (round_Signal[1]), .Z0_t (Midori_rounds_constant_MUX_n69) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U5 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n34), .Z0_t (Midori_rounds_constant_MUX_n50) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U4 ( .A0_t (enc_dec), .B0_t (round_Signal[0]), .Z0_t (Midori_rounds_constant_MUX_n34) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U2 ( .A0_t (round_Signal[2]), .B0_t (Midori_rounds_constant_MUX_n56), .Z0_t (Midori_rounds_constant_MUX_n111) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U1 ( .A0_t (round_Signal[0]), .B0_t (enc_dec), .Z0_t (Midori_rounds_constant_MUX_n56) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U53_XOR1_U1 ( .A0_t (Midori_rounds_constant_MUX_n121), .B0_t (Midori_rounds_constant_MUX_n111), .Z0_t (Midori_rounds_constant_MUX_U53_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U53_AND1_U1 ( .A0_t (round_Signal[3]), .B0_t (Midori_rounds_constant_MUX_U53_X), .Z0_t (Midori_rounds_constant_MUX_U53_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U53_XOR2_U1 ( .A0_t (Midori_rounds_constant_MUX_U53_Y), .B0_t (Midori_rounds_constant_MUX_n121), .Z0_t (Midori_rounds_constant_MUX_n43) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U119_XOR1_U1 ( .A0_t (Midori_rounds_constant_MUX_n111), .B0_t (Midori_rounds_constant_MUX_n121), .Z0_t (Midori_rounds_constant_MUX_U119_X) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b1)) Midori_rounds_constant_MUX_U119_AND1_U1 ( .A0_t (round_Signal[3]), .B0_t (Midori_rounds_constant_MUX_U119_X), .Z0_t (Midori_rounds_constant_MUX_U119_Y) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0), .NL(1'b0)) Midori_rounds_constant_MUX_U119_XOR2_U1 ( .A0_t (Midori_rounds_constant_MUX_U119_Y), .B0_t (Midori_rounds_constant_MUX_n111), .Z0_t (Midori_rounds_constant_MUX_n112) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_XOR1_U1 ( .A0_t (key[64]), .B0_t (key[0]), .Z0_t (Midori_rounds_MUXInst_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_0_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_0_U1_Y), .B0_t (key[64]), .Z0_t (Midori_rounds_SelectedKey[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_XOR1_U1 ( .A0_t (key[65]), .B0_t (key[1]), .Z0_t (Midori_rounds_MUXInst_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_1_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_1_U1_Y), .B0_t (key[65]), .Z0_t (Midori_rounds_SelectedKey[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_XOR1_U1 ( .A0_t (key[66]), .B0_t (key[2]), .Z0_t (Midori_rounds_MUXInst_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_2_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_2_U1_Y), .B0_t (key[66]), .Z0_t (Midori_rounds_SelectedKey[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_XOR1_U1 ( .A0_t (key[67]), .B0_t (key[3]), .Z0_t (Midori_rounds_MUXInst_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_3_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_3_U1_Y), .B0_t (key[67]), .Z0_t (Midori_rounds_SelectedKey[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_XOR1_U1 ( .A0_t (key[68]), .B0_t (key[4]), .Z0_t (Midori_rounds_MUXInst_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_4_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_4_U1_Y), .B0_t (key[68]), .Z0_t (Midori_rounds_SelectedKey[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_XOR1_U1 ( .A0_t (key[69]), .B0_t (key[5]), .Z0_t (Midori_rounds_MUXInst_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_5_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_5_U1_Y), .B0_t (key[69]), .Z0_t (Midori_rounds_SelectedKey[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_XOR1_U1 ( .A0_t (key[70]), .B0_t (key[6]), .Z0_t (Midori_rounds_MUXInst_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_6_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_6_U1_Y), .B0_t (key[70]), .Z0_t (Midori_rounds_SelectedKey[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_XOR1_U1 ( .A0_t (key[71]), .B0_t (key[7]), .Z0_t (Midori_rounds_MUXInst_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_7_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_7_U1_Y), .B0_t (key[71]), .Z0_t (Midori_rounds_SelectedKey[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_XOR1_U1 ( .A0_t (key[72]), .B0_t (key[8]), .Z0_t (Midori_rounds_MUXInst_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_8_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_8_U1_Y), .B0_t (key[72]), .Z0_t (Midori_rounds_SelectedKey[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_XOR1_U1 ( .A0_t (key[73]), .B0_t (key[9]), .Z0_t (Midori_rounds_MUXInst_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_9_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_9_U1_Y), .B0_t (key[73]), .Z0_t (Midori_rounds_SelectedKey[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_XOR1_U1 ( .A0_t (key[74]), .B0_t (key[10]), .Z0_t (Midori_rounds_MUXInst_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_10_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_10_U1_Y), .B0_t (key[74]), .Z0_t (Midori_rounds_SelectedKey[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_XOR1_U1 ( .A0_t (key[75]), .B0_t (key[11]), .Z0_t (Midori_rounds_MUXInst_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_11_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_11_U1_Y), .B0_t (key[75]), .Z0_t (Midori_rounds_SelectedKey[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_XOR1_U1 ( .A0_t (key[76]), .B0_t (key[12]), .Z0_t (Midori_rounds_MUXInst_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_12_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_12_U1_Y), .B0_t (key[76]), .Z0_t (Midori_rounds_SelectedKey[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_XOR1_U1 ( .A0_t (key[77]), .B0_t (key[13]), .Z0_t (Midori_rounds_MUXInst_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_13_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_13_U1_Y), .B0_t (key[77]), .Z0_t (Midori_rounds_SelectedKey[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_XOR1_U1 ( .A0_t (key[78]), .B0_t (key[14]), .Z0_t (Midori_rounds_MUXInst_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_14_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_14_U1_Y), .B0_t (key[78]), .Z0_t (Midori_rounds_SelectedKey[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_XOR1_U1 ( .A0_t (key[79]), .B0_t (key[15]), .Z0_t (Midori_rounds_MUXInst_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_15_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_15_U1_Y), .B0_t (key[79]), .Z0_t (Midori_rounds_SelectedKey[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_XOR1_U1 ( .A0_t (key[80]), .B0_t (key[16]), .Z0_t (Midori_rounds_MUXInst_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_16_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_16_U1_Y), .B0_t (key[80]), .Z0_t (Midori_rounds_SelectedKey[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_XOR1_U1 ( .A0_t (key[81]), .B0_t (key[17]), .Z0_t (Midori_rounds_MUXInst_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_17_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_17_U1_Y), .B0_t (key[81]), .Z0_t (Midori_rounds_SelectedKey[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_XOR1_U1 ( .A0_t (key[82]), .B0_t (key[18]), .Z0_t (Midori_rounds_MUXInst_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_18_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_18_U1_Y), .B0_t (key[82]), .Z0_t (Midori_rounds_SelectedKey[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_XOR1_U1 ( .A0_t (key[83]), .B0_t (key[19]), .Z0_t (Midori_rounds_MUXInst_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_19_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_19_U1_Y), .B0_t (key[83]), .Z0_t (Midori_rounds_SelectedKey[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_XOR1_U1 ( .A0_t (key[84]), .B0_t (key[20]), .Z0_t (Midori_rounds_MUXInst_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_20_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_20_U1_Y), .B0_t (key[84]), .Z0_t (Midori_rounds_SelectedKey[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_XOR1_U1 ( .A0_t (key[85]), .B0_t (key[21]), .Z0_t (Midori_rounds_MUXInst_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_21_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_21_U1_Y), .B0_t (key[85]), .Z0_t (Midori_rounds_SelectedKey[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_XOR1_U1 ( .A0_t (key[86]), .B0_t (key[22]), .Z0_t (Midori_rounds_MUXInst_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_22_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_22_U1_Y), .B0_t (key[86]), .Z0_t (Midori_rounds_SelectedKey[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_XOR1_U1 ( .A0_t (key[87]), .B0_t (key[23]), .Z0_t (Midori_rounds_MUXInst_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_23_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_23_U1_Y), .B0_t (key[87]), .Z0_t (Midori_rounds_SelectedKey[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_XOR1_U1 ( .A0_t (key[88]), .B0_t (key[24]), .Z0_t (Midori_rounds_MUXInst_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_24_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_24_U1_Y), .B0_t (key[88]), .Z0_t (Midori_rounds_SelectedKey[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_XOR1_U1 ( .A0_t (key[89]), .B0_t (key[25]), .Z0_t (Midori_rounds_MUXInst_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_25_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_25_U1_Y), .B0_t (key[89]), .Z0_t (Midori_rounds_SelectedKey[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_XOR1_U1 ( .A0_t (key[90]), .B0_t (key[26]), .Z0_t (Midori_rounds_MUXInst_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_26_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_26_U1_Y), .B0_t (key[90]), .Z0_t (Midori_rounds_SelectedKey[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_XOR1_U1 ( .A0_t (key[91]), .B0_t (key[27]), .Z0_t (Midori_rounds_MUXInst_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_27_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_27_U1_Y), .B0_t (key[91]), .Z0_t (Midori_rounds_SelectedKey[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_XOR1_U1 ( .A0_t (key[92]), .B0_t (key[28]), .Z0_t (Midori_rounds_MUXInst_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_28_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_28_U1_Y), .B0_t (key[92]), .Z0_t (Midori_rounds_SelectedKey[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_XOR1_U1 ( .A0_t (key[93]), .B0_t (key[29]), .Z0_t (Midori_rounds_MUXInst_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_29_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_29_U1_Y), .B0_t (key[93]), .Z0_t (Midori_rounds_SelectedKey[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_XOR1_U1 ( .A0_t (key[94]), .B0_t (key[30]), .Z0_t (Midori_rounds_MUXInst_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_30_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_30_U1_Y), .B0_t (key[94]), .Z0_t (Midori_rounds_SelectedKey[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_XOR1_U1 ( .A0_t (key[95]), .B0_t (key[31]), .Z0_t (Midori_rounds_MUXInst_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_31_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_31_U1_Y), .B0_t (key[95]), .Z0_t (Midori_rounds_SelectedKey[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_XOR1_U1 ( .A0_t (key[96]), .B0_t (key[32]), .Z0_t (Midori_rounds_MUXInst_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_32_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_32_U1_Y), .B0_t (key[96]), .Z0_t (Midori_rounds_SelectedKey[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_XOR1_U1 ( .A0_t (key[97]), .B0_t (key[33]), .Z0_t (Midori_rounds_MUXInst_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_33_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_33_U1_Y), .B0_t (key[97]), .Z0_t (Midori_rounds_SelectedKey[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_XOR1_U1 ( .A0_t (key[98]), .B0_t (key[34]), .Z0_t (Midori_rounds_MUXInst_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_34_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_34_U1_Y), .B0_t (key[98]), .Z0_t (Midori_rounds_SelectedKey[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_XOR1_U1 ( .A0_t (key[99]), .B0_t (key[35]), .Z0_t (Midori_rounds_MUXInst_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_35_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_35_U1_Y), .B0_t (key[99]), .Z0_t (Midori_rounds_SelectedKey[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_XOR1_U1 ( .A0_t (key[100]), .B0_t (key[36]), .Z0_t (Midori_rounds_MUXInst_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_36_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_36_U1_Y), .B0_t (key[100]), .Z0_t (Midori_rounds_SelectedKey[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_XOR1_U1 ( .A0_t (key[101]), .B0_t (key[37]), .Z0_t (Midori_rounds_MUXInst_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_37_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_37_U1_Y), .B0_t (key[101]), .Z0_t (Midori_rounds_SelectedKey[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_XOR1_U1 ( .A0_t (key[102]), .B0_t (key[38]), .Z0_t (Midori_rounds_MUXInst_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_38_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_38_U1_Y), .B0_t (key[102]), .Z0_t (Midori_rounds_SelectedKey[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_XOR1_U1 ( .A0_t (key[103]), .B0_t (key[39]), .Z0_t (Midori_rounds_MUXInst_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_39_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_39_U1_Y), .B0_t (key[103]), .Z0_t (Midori_rounds_SelectedKey[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_XOR1_U1 ( .A0_t (key[104]), .B0_t (key[40]), .Z0_t (Midori_rounds_MUXInst_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_40_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_40_U1_Y), .B0_t (key[104]), .Z0_t (Midori_rounds_SelectedKey[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_XOR1_U1 ( .A0_t (key[105]), .B0_t (key[41]), .Z0_t (Midori_rounds_MUXInst_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_41_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_41_U1_Y), .B0_t (key[105]), .Z0_t (Midori_rounds_SelectedKey[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_XOR1_U1 ( .A0_t (key[106]), .B0_t (key[42]), .Z0_t (Midori_rounds_MUXInst_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_42_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_42_U1_Y), .B0_t (key[106]), .Z0_t (Midori_rounds_SelectedKey[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_XOR1_U1 ( .A0_t (key[107]), .B0_t (key[43]), .Z0_t (Midori_rounds_MUXInst_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_43_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_43_U1_Y), .B0_t (key[107]), .Z0_t (Midori_rounds_SelectedKey[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_XOR1_U1 ( .A0_t (key[108]), .B0_t (key[44]), .Z0_t (Midori_rounds_MUXInst_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_44_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_44_U1_Y), .B0_t (key[108]), .Z0_t (Midori_rounds_SelectedKey[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_XOR1_U1 ( .A0_t (key[109]), .B0_t (key[45]), .Z0_t (Midori_rounds_MUXInst_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_45_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_45_U1_Y), .B0_t (key[109]), .Z0_t (Midori_rounds_SelectedKey[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_XOR1_U1 ( .A0_t (key[110]), .B0_t (key[46]), .Z0_t (Midori_rounds_MUXInst_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_46_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_46_U1_Y), .B0_t (key[110]), .Z0_t (Midori_rounds_SelectedKey[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_XOR1_U1 ( .A0_t (key[111]), .B0_t (key[47]), .Z0_t (Midori_rounds_MUXInst_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_47_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_47_U1_Y), .B0_t (key[111]), .Z0_t (Midori_rounds_SelectedKey[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_XOR1_U1 ( .A0_t (key[112]), .B0_t (key[48]), .Z0_t (Midori_rounds_MUXInst_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_48_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_48_U1_Y), .B0_t (key[112]), .Z0_t (Midori_rounds_SelectedKey[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_XOR1_U1 ( .A0_t (key[113]), .B0_t (key[49]), .Z0_t (Midori_rounds_MUXInst_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_49_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_49_U1_Y), .B0_t (key[113]), .Z0_t (Midori_rounds_SelectedKey[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_XOR1_U1 ( .A0_t (key[114]), .B0_t (key[50]), .Z0_t (Midori_rounds_MUXInst_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_50_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_50_U1_Y), .B0_t (key[114]), .Z0_t (Midori_rounds_SelectedKey[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_XOR1_U1 ( .A0_t (key[115]), .B0_t (key[51]), .Z0_t (Midori_rounds_MUXInst_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_51_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_51_U1_Y), .B0_t (key[115]), .Z0_t (Midori_rounds_SelectedKey[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_XOR1_U1 ( .A0_t (key[116]), .B0_t (key[52]), .Z0_t (Midori_rounds_MUXInst_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_52_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_52_U1_Y), .B0_t (key[116]), .Z0_t (Midori_rounds_SelectedKey[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_XOR1_U1 ( .A0_t (key[117]), .B0_t (key[53]), .Z0_t (Midori_rounds_MUXInst_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_53_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_53_U1_Y), .B0_t (key[117]), .Z0_t (Midori_rounds_SelectedKey[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_XOR1_U1 ( .A0_t (key[118]), .B0_t (key[54]), .Z0_t (Midori_rounds_MUXInst_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_54_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_54_U1_Y), .B0_t (key[118]), .Z0_t (Midori_rounds_SelectedKey[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_XOR1_U1 ( .A0_t (key[119]), .B0_t (key[55]), .Z0_t (Midori_rounds_MUXInst_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_55_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_55_U1_Y), .B0_t (key[119]), .Z0_t (Midori_rounds_SelectedKey[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_XOR1_U1 ( .A0_t (key[120]), .B0_t (key[56]), .Z0_t (Midori_rounds_MUXInst_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_56_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_56_U1_Y), .B0_t (key[120]), .Z0_t (Midori_rounds_SelectedKey[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_XOR1_U1 ( .A0_t (key[121]), .B0_t (key[57]), .Z0_t (Midori_rounds_MUXInst_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_57_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_57_U1_Y), .B0_t (key[121]), .Z0_t (Midori_rounds_SelectedKey[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_XOR1_U1 ( .A0_t (key[122]), .B0_t (key[58]), .Z0_t (Midori_rounds_MUXInst_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_58_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_58_U1_Y), .B0_t (key[122]), .Z0_t (Midori_rounds_SelectedKey[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_XOR1_U1 ( .A0_t (key[123]), .B0_t (key[59]), .Z0_t (Midori_rounds_MUXInst_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_59_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_59_U1_Y), .B0_t (key[123]), .Z0_t (Midori_rounds_SelectedKey[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_XOR1_U1 ( .A0_t (key[124]), .B0_t (key[60]), .Z0_t (Midori_rounds_MUXInst_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_60_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_60_U1_Y), .B0_t (key[124]), .Z0_t (Midori_rounds_SelectedKey[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_XOR1_U1 ( .A0_t (key[125]), .B0_t (key[61]), .Z0_t (Midori_rounds_MUXInst_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_61_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_61_U1_Y), .B0_t (key[125]), .Z0_t (Midori_rounds_SelectedKey[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_XOR1_U1 ( .A0_t (key[126]), .B0_t (key[62]), .Z0_t (Midori_rounds_MUXInst_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_62_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_62_U1_Y), .B0_t (key[126]), .Z0_t (Midori_rounds_SelectedKey[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_XOR1_U1 ( .A0_t (key[127]), .B0_t (key[63]), .Z0_t (Midori_rounds_MUXInst_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_AND1_U1 ( .A0_t (round_Signal[0]), .B0_t (Midori_rounds_MUXInst_mux_inst_63_U1_X), .Z0_t (Midori_rounds_MUXInst_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_MUXInst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_MUXInst_mux_inst_63_U1_Y), .B0_t (key[127]), .Z0_t (Midori_rounds_SelectedKey[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[0]), .B0_t (Midori_add_Result_Start[0]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_0_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[0]), .Z0_t (Midori_rounds_roundReg_out[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[1]), .B0_t (Midori_add_Result_Start[1]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_1_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[1]), .Z0_t (Midori_rounds_roundReg_out[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[2]), .B0_t (Midori_add_Result_Start[2]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_2_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[2]), .Z0_t (Midori_rounds_roundReg_out[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[3]), .B0_t (Midori_add_Result_Start[3]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_3_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[3]), .Z0_t (Midori_rounds_roundReg_out[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[4]), .B0_t (Midori_add_Result_Start[4]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_4_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[4]), .Z0_t (Midori_rounds_roundReg_out[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[5]), .B0_t (Midori_add_Result_Start[5]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_5_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[5]), .Z0_t (Midori_rounds_roundReg_out[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[6]), .B0_t (Midori_add_Result_Start[6]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_6_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[6]), .Z0_t (Midori_rounds_roundReg_out[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[7]), .B0_t (Midori_add_Result_Start[7]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_7_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[7]), .Z0_t (Midori_rounds_roundReg_out[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[8]), .B0_t (Midori_add_Result_Start[8]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_8_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[8]), .Z0_t (Midori_rounds_roundReg_out[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[9]), .B0_t (Midori_add_Result_Start[9]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_9_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[9]), .Z0_t (Midori_rounds_roundReg_out[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[10]), .B0_t (Midori_add_Result_Start[10]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_10_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[10]), .Z0_t (Midori_rounds_roundReg_out[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[11]), .B0_t (Midori_add_Result_Start[11]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_11_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[11]), .Z0_t (Midori_rounds_roundReg_out[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[12]), .B0_t (Midori_add_Result_Start[12]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_12_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[12]), .Z0_t (Midori_rounds_roundReg_out[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[13]), .B0_t (Midori_add_Result_Start[13]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_13_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[13]), .Z0_t (Midori_rounds_roundReg_out[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[14]), .B0_t (Midori_add_Result_Start[14]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_14_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[14]), .Z0_t (Midori_rounds_roundReg_out[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[15]), .B0_t (Midori_add_Result_Start[15]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_15_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[15]), .Z0_t (Midori_rounds_roundReg_out[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[16]), .B0_t (Midori_add_Result_Start[16]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_16_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[16]), .Z0_t (Midori_rounds_roundReg_out[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[17]), .B0_t (Midori_add_Result_Start[17]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_17_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[17]), .Z0_t (Midori_rounds_roundReg_out[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[18]), .B0_t (Midori_add_Result_Start[18]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_18_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[18]), .Z0_t (Midori_rounds_roundReg_out[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[19]), .B0_t (Midori_add_Result_Start[19]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_19_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[19]), .Z0_t (Midori_rounds_roundReg_out[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[20]), .B0_t (Midori_add_Result_Start[20]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_20_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[20]), .Z0_t (Midori_rounds_roundReg_out[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[21]), .B0_t (Midori_add_Result_Start[21]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_21_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[21]), .Z0_t (Midori_rounds_roundReg_out[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[22]), .B0_t (Midori_add_Result_Start[22]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_22_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[22]), .Z0_t (Midori_rounds_roundReg_out[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[23]), .B0_t (Midori_add_Result_Start[23]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_23_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[23]), .Z0_t (Midori_rounds_roundReg_out[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[24]), .B0_t (Midori_add_Result_Start[24]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_24_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[24]), .Z0_t (Midori_rounds_roundReg_out[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[25]), .B0_t (Midori_add_Result_Start[25]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_25_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[25]), .Z0_t (Midori_rounds_roundReg_out[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[26]), .B0_t (Midori_add_Result_Start[26]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_26_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[26]), .Z0_t (Midori_rounds_roundReg_out[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[27]), .B0_t (Midori_add_Result_Start[27]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_27_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[27]), .Z0_t (Midori_rounds_roundReg_out[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[28]), .B0_t (Midori_add_Result_Start[28]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_28_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[28]), .Z0_t (Midori_rounds_roundReg_out[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[29]), .B0_t (Midori_add_Result_Start[29]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_29_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[29]), .Z0_t (Midori_rounds_roundReg_out[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[30]), .B0_t (Midori_add_Result_Start[30]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_30_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[30]), .Z0_t (Midori_rounds_roundReg_out[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[31]), .B0_t (Midori_add_Result_Start[31]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_31_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[31]), .Z0_t (Midori_rounds_roundReg_out[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[32]), .B0_t (Midori_add_Result_Start[32]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_32_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[32]), .Z0_t (Midori_rounds_roundReg_out[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[33]), .B0_t (Midori_add_Result_Start[33]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_33_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[33]), .Z0_t (Midori_rounds_roundReg_out[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[34]), .B0_t (Midori_add_Result_Start[34]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_34_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[34]), .Z0_t (Midori_rounds_roundReg_out[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[35]), .B0_t (Midori_add_Result_Start[35]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_35_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[35]), .Z0_t (Midori_rounds_roundReg_out[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[36]), .B0_t (Midori_add_Result_Start[36]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_36_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[36]), .Z0_t (Midori_rounds_roundReg_out[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[37]), .B0_t (Midori_add_Result_Start[37]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_37_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[37]), .Z0_t (Midori_rounds_roundReg_out[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[38]), .B0_t (Midori_add_Result_Start[38]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_38_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[38]), .Z0_t (Midori_rounds_roundReg_out[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[39]), .B0_t (Midori_add_Result_Start[39]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_39_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[39]), .Z0_t (Midori_rounds_roundReg_out[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[40]), .B0_t (Midori_add_Result_Start[40]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_40_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[40]), .Z0_t (Midori_rounds_roundReg_out[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[41]), .B0_t (Midori_add_Result_Start[41]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_41_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[41]), .Z0_t (Midori_rounds_roundReg_out[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[42]), .B0_t (Midori_add_Result_Start[42]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_42_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[42]), .Z0_t (Midori_rounds_roundReg_out[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[43]), .B0_t (Midori_add_Result_Start[43]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_43_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[43]), .Z0_t (Midori_rounds_roundReg_out[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[44]), .B0_t (Midori_add_Result_Start[44]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_44_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[44]), .Z0_t (Midori_rounds_roundReg_out[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[45]), .B0_t (Midori_add_Result_Start[45]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_45_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[45]), .Z0_t (Midori_rounds_roundReg_out[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[46]), .B0_t (Midori_add_Result_Start[46]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_46_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[46]), .Z0_t (Midori_rounds_roundReg_out[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[47]), .B0_t (Midori_add_Result_Start[47]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_47_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[47]), .Z0_t (Midori_rounds_roundReg_out[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[48]), .B0_t (Midori_add_Result_Start[48]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_48_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[48]), .Z0_t (Midori_rounds_roundReg_out[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[49]), .B0_t (Midori_add_Result_Start[49]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_49_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[49]), .Z0_t (Midori_rounds_roundReg_out[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[50]), .B0_t (Midori_add_Result_Start[50]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_50_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[50]), .Z0_t (Midori_rounds_roundReg_out[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[51]), .B0_t (Midori_add_Result_Start[51]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_51_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[51]), .Z0_t (Midori_rounds_roundReg_out[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[52]), .B0_t (Midori_add_Result_Start[52]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_52_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[52]), .Z0_t (Midori_rounds_roundReg_out[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[53]), .B0_t (Midori_add_Result_Start[53]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_53_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[53]), .Z0_t (Midori_rounds_roundReg_out[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[54]), .B0_t (Midori_add_Result_Start[54]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_54_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[54]), .Z0_t (Midori_rounds_roundReg_out[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[55]), .B0_t (Midori_add_Result_Start[55]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_55_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[55]), .Z0_t (Midori_rounds_roundReg_out[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[56]), .B0_t (Midori_add_Result_Start[56]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_56_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[56]), .Z0_t (Midori_rounds_roundReg_out[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[57]), .B0_t (Midori_add_Result_Start[57]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_57_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[57]), .Z0_t (Midori_rounds_roundReg_out[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[58]), .B0_t (Midori_add_Result_Start[58]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_58_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[58]), .Z0_t (Midori_rounds_roundReg_out[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[59]), .B0_t (Midori_add_Result_Start[59]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_59_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[59]), .Z0_t (Midori_rounds_roundReg_out[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[60]), .B0_t (Midori_add_Result_Start[60]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_60_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[60]), .Z0_t (Midori_rounds_roundReg_out[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[61]), .B0_t (Midori_add_Result_Start[61]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_61_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[61]), .Z0_t (Midori_rounds_roundReg_out[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[62]), .B0_t (Midori_add_Result_Start[62]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_62_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[62]), .Z0_t (Midori_rounds_roundReg_out[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_XOR1_U1 ( .A0_t (Midori_rounds_round_Result[63]), .B0_t (Midori_add_Result_Start[63]), .Z0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_AND1_U1 ( .A0_t (reset), .B0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_X), .Z0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1)) Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_XOR2_U1 ( .A0_t (Midori_rounds_roundResult_Reg_SFF_63_MUXInst_U1_Y), .B0_t (Midori_rounds_round_Result[63]), .Z0_t (Midori_rounds_roundReg_out[63]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n14), .Z0_t (Midori_rounds_SR_Result[51]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n13), .B0_t (Midori_rounds_roundReg_out[1]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n11), .Z0_t (Midori_rounds_SR_Result[49]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U16 ( .A0_t (Midori_rounds_roundReg_out[0]), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U15 ( .A0_t (Midori_rounds_roundReg_out[3]), .B0_t (Midori_rounds_roundReg_out[2]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U14 ( .A0_t (Midori_rounds_roundReg_out[2]), .B0_t (Midori_rounds_roundReg_out[3]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n7), .Z0_t (Midori_rounds_SR_Result[50]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n6), .B0_t (Midori_rounds_roundReg_out[1]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n5), .B0_t (Midori_rounds_roundReg_out[2]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U10 ( .A0_t (Midori_rounds_roundReg_out[0]), .B0_t (Midori_rounds_roundReg_out[3]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U9 ( .A0_t (Midori_rounds_roundReg_out[3]), .B0_t (Midori_rounds_roundReg_out[0]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_0_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n3), .Z0_t (Midori_rounds_SR_Result[48]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U7 ( .A0_t (Midori_rounds_roundReg_out[1]), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U6 ( .A0_t (Midori_rounds_roundReg_out[0]), .B0_t (Midori_rounds_sub_sBox_PRINCE_0_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U5 ( .A0_t (Midori_rounds_roundReg_out[2]), .B0_t (Midori_rounds_roundReg_out[3]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_0_U3 ( .A0_t (Midori_rounds_roundReg_out[2]), .B0_t (Midori_rounds_roundReg_out[3]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_0_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n14), .Z0_t (Midori_rounds_SR_Result[44]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U18 ( .A0_t (Midori_rounds_roundReg_out[5]), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U17 ( .A0_t (Midori_rounds_roundReg_out[4]), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U16 ( .A0_t (Midori_rounds_roundReg_out[6]), .B0_t (Midori_rounds_roundReg_out[7]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n9), .Z0_t (Midori_rounds_SR_Result[46]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n8), .B0_t (Midori_rounds_roundReg_out[5]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n7), .B0_t (Midori_rounds_roundReg_out[6]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U12 ( .A0_t (Midori_rounds_roundReg_out[4]), .B0_t (Midori_rounds_roundReg_out[7]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n5), .Z0_t (Midori_rounds_SR_Result[47]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U10 ( .A0_t (Midori_rounds_roundReg_out[5]), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U9 ( .A0_t (Midori_rounds_roundReg_out[6]), .B0_t (Midori_rounds_roundReg_out[7]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U8 ( .A0_t (Midori_rounds_roundReg_out[7]), .B0_t (Midori_rounds_roundReg_out[4]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_1_n2), .Z0_t (Midori_rounds_SR_Result[45]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_1_n1), .B0_t (Midori_rounds_roundReg_out[7]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U4 ( .A0_t (Midori_rounds_roundReg_out[6]), .B0_t (Midori_rounds_roundReg_out[4]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_1_U1 ( .A0_t (Midori_rounds_roundReg_out[6]), .B0_t (Midori_rounds_roundReg_out[4]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_1_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n14), .Z0_t (Midori_rounds_SR_Result[8]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U18 ( .A0_t (Midori_rounds_roundReg_out[9]), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U17 ( .A0_t (Midori_rounds_roundReg_out[8]), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U16 ( .A0_t (Midori_rounds_roundReg_out[10]), .B0_t (Midori_rounds_roundReg_out[11]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n9), .Z0_t (Midori_rounds_SR_Result[10]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n8), .B0_t (Midori_rounds_roundReg_out[9]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n7), .B0_t (Midori_rounds_roundReg_out[10]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U12 ( .A0_t (Midori_rounds_roundReg_out[8]), .B0_t (Midori_rounds_roundReg_out[11]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n5), .Z0_t (Midori_rounds_SR_Result[11]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U10 ( .A0_t (Midori_rounds_roundReg_out[9]), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U9 ( .A0_t (Midori_rounds_roundReg_out[10]), .B0_t (Midori_rounds_roundReg_out[11]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U8 ( .A0_t (Midori_rounds_roundReg_out[11]), .B0_t (Midori_rounds_roundReg_out[8]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_2_n2), .Z0_t (Midori_rounds_SR_Result[9]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_2_n1), .B0_t (Midori_rounds_roundReg_out[11]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U4 ( .A0_t (Midori_rounds_roundReg_out[10]), .B0_t (Midori_rounds_roundReg_out[8]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_2_U1 ( .A0_t (Midori_rounds_roundReg_out[10]), .B0_t (Midori_rounds_roundReg_out[8]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_2_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n14), .Z0_t (Midori_rounds_SR_Result[20]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U18 ( .A0_t (Midori_rounds_roundReg_out[13]), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U17 ( .A0_t (Midori_rounds_roundReg_out[12]), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U16 ( .A0_t (Midori_rounds_roundReg_out[14]), .B0_t (Midori_rounds_roundReg_out[15]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n9), .Z0_t (Midori_rounds_SR_Result[22]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n8), .B0_t (Midori_rounds_roundReg_out[13]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n7), .B0_t (Midori_rounds_roundReg_out[14]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U12 ( .A0_t (Midori_rounds_roundReg_out[12]), .B0_t (Midori_rounds_roundReg_out[15]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n5), .Z0_t (Midori_rounds_SR_Result[23]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U10 ( .A0_t (Midori_rounds_roundReg_out[13]), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U9 ( .A0_t (Midori_rounds_roundReg_out[14]), .B0_t (Midori_rounds_roundReg_out[15]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U8 ( .A0_t (Midori_rounds_roundReg_out[15]), .B0_t (Midori_rounds_roundReg_out[12]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_3_n2), .Z0_t (Midori_rounds_SR_Result[21]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_3_n1), .B0_t (Midori_rounds_roundReg_out[15]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U4 ( .A0_t (Midori_rounds_roundReg_out[14]), .B0_t (Midori_rounds_roundReg_out[12]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_3_U1 ( .A0_t (Midori_rounds_roundReg_out[14]), .B0_t (Midori_rounds_roundReg_out[12]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_3_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n14), .Z0_t (Midori_rounds_SR_Result[36]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U18 ( .A0_t (Midori_rounds_roundReg_out[17]), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U17 ( .A0_t (Midori_rounds_roundReg_out[16]), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U16 ( .A0_t (Midori_rounds_roundReg_out[18]), .B0_t (Midori_rounds_roundReg_out[19]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n9), .Z0_t (Midori_rounds_SR_Result[38]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n8), .B0_t (Midori_rounds_roundReg_out[17]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n7), .B0_t (Midori_rounds_roundReg_out[18]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U12 ( .A0_t (Midori_rounds_roundReg_out[16]), .B0_t (Midori_rounds_roundReg_out[19]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n5), .Z0_t (Midori_rounds_SR_Result[39]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U10 ( .A0_t (Midori_rounds_roundReg_out[17]), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U9 ( .A0_t (Midori_rounds_roundReg_out[18]), .B0_t (Midori_rounds_roundReg_out[19]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U8 ( .A0_t (Midori_rounds_roundReg_out[19]), .B0_t (Midori_rounds_roundReg_out[16]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_4_n2), .Z0_t (Midori_rounds_SR_Result[37]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_4_n1), .B0_t (Midori_rounds_roundReg_out[19]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U4 ( .A0_t (Midori_rounds_roundReg_out[18]), .B0_t (Midori_rounds_roundReg_out[16]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_4_U1 ( .A0_t (Midori_rounds_roundReg_out[18]), .B0_t (Midori_rounds_roundReg_out[16]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_4_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n14), .Z0_t (Midori_rounds_SR_Result[56]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U18 ( .A0_t (Midori_rounds_roundReg_out[21]), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U17 ( .A0_t (Midori_rounds_roundReg_out[20]), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U16 ( .A0_t (Midori_rounds_roundReg_out[22]), .B0_t (Midori_rounds_roundReg_out[23]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n9), .Z0_t (Midori_rounds_SR_Result[58]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n8), .B0_t (Midori_rounds_roundReg_out[21]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n7), .B0_t (Midori_rounds_roundReg_out[22]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U12 ( .A0_t (Midori_rounds_roundReg_out[20]), .B0_t (Midori_rounds_roundReg_out[23]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n5), .Z0_t (Midori_rounds_SR_Result[59]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U10 ( .A0_t (Midori_rounds_roundReg_out[21]), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U9 ( .A0_t (Midori_rounds_roundReg_out[22]), .B0_t (Midori_rounds_roundReg_out[23]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U8 ( .A0_t (Midori_rounds_roundReg_out[23]), .B0_t (Midori_rounds_roundReg_out[20]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_5_n2), .Z0_t (Midori_rounds_SR_Result[57]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_5_n1), .B0_t (Midori_rounds_roundReg_out[23]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U4 ( .A0_t (Midori_rounds_roundReg_out[22]), .B0_t (Midori_rounds_roundReg_out[20]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_5_U1 ( .A0_t (Midori_rounds_roundReg_out[22]), .B0_t (Midori_rounds_roundReg_out[20]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_5_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n14), .Z0_t (Midori_rounds_SR_Result[28]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U18 ( .A0_t (Midori_rounds_roundReg_out[25]), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U17 ( .A0_t (Midori_rounds_roundReg_out[24]), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U16 ( .A0_t (Midori_rounds_roundReg_out[26]), .B0_t (Midori_rounds_roundReg_out[27]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n9), .Z0_t (Midori_rounds_SR_Result[30]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n8), .B0_t (Midori_rounds_roundReg_out[25]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n7), .B0_t (Midori_rounds_roundReg_out[26]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U12 ( .A0_t (Midori_rounds_roundReg_out[24]), .B0_t (Midori_rounds_roundReg_out[27]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n5), .Z0_t (Midori_rounds_SR_Result[31]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U10 ( .A0_t (Midori_rounds_roundReg_out[25]), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U9 ( .A0_t (Midori_rounds_roundReg_out[26]), .B0_t (Midori_rounds_roundReg_out[27]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U8 ( .A0_t (Midori_rounds_roundReg_out[27]), .B0_t (Midori_rounds_roundReg_out[24]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_6_n2), .Z0_t (Midori_rounds_SR_Result[29]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_6_n1), .B0_t (Midori_rounds_roundReg_out[27]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U4 ( .A0_t (Midori_rounds_roundReg_out[26]), .B0_t (Midori_rounds_roundReg_out[24]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_6_U1 ( .A0_t (Midori_rounds_roundReg_out[26]), .B0_t (Midori_rounds_roundReg_out[24]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_6_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n14), .Z0_t (Midori_rounds_SR_Result[3]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n13), .B0_t (Midori_rounds_roundReg_out[29]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n11), .Z0_t (Midori_rounds_SR_Result[1]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U16 ( .A0_t (Midori_rounds_roundReg_out[28]), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U15 ( .A0_t (Midori_rounds_roundReg_out[31]), .B0_t (Midori_rounds_roundReg_out[30]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U14 ( .A0_t (Midori_rounds_roundReg_out[30]), .B0_t (Midori_rounds_roundReg_out[31]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n7), .Z0_t (Midori_rounds_SR_Result[2]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n6), .B0_t (Midori_rounds_roundReg_out[29]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n5), .B0_t (Midori_rounds_roundReg_out[30]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U10 ( .A0_t (Midori_rounds_roundReg_out[28]), .B0_t (Midori_rounds_roundReg_out[31]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U9 ( .A0_t (Midori_rounds_roundReg_out[31]), .B0_t (Midori_rounds_roundReg_out[28]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_7_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n3), .Z0_t (Midori_rounds_SR_Result[0]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U7 ( .A0_t (Midori_rounds_roundReg_out[29]), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U6 ( .A0_t (Midori_rounds_roundReg_out[28]), .B0_t (Midori_rounds_sub_sBox_PRINCE_7_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U5 ( .A0_t (Midori_rounds_roundReg_out[30]), .B0_t (Midori_rounds_roundReg_out[31]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_7_U3 ( .A0_t (Midori_rounds_roundReg_out[30]), .B0_t (Midori_rounds_roundReg_out[31]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_7_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n14), .Z0_t (Midori_rounds_SR_Result[15]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n13), .B0_t (Midori_rounds_roundReg_out[33]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n11), .Z0_t (Midori_rounds_SR_Result[13]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U16 ( .A0_t (Midori_rounds_roundReg_out[32]), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U15 ( .A0_t (Midori_rounds_roundReg_out[35]), .B0_t (Midori_rounds_roundReg_out[34]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U14 ( .A0_t (Midori_rounds_roundReg_out[34]), .B0_t (Midori_rounds_roundReg_out[35]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n7), .Z0_t (Midori_rounds_SR_Result[14]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n6), .B0_t (Midori_rounds_roundReg_out[33]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n5), .B0_t (Midori_rounds_roundReg_out[34]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U10 ( .A0_t (Midori_rounds_roundReg_out[32]), .B0_t (Midori_rounds_roundReg_out[35]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U9 ( .A0_t (Midori_rounds_roundReg_out[35]), .B0_t (Midori_rounds_roundReg_out[32]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_8_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n3), .Z0_t (Midori_rounds_SR_Result[12]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U7 ( .A0_t (Midori_rounds_roundReg_out[33]), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U6 ( .A0_t (Midori_rounds_roundReg_out[32]), .B0_t (Midori_rounds_sub_sBox_PRINCE_8_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U5 ( .A0_t (Midori_rounds_roundReg_out[34]), .B0_t (Midori_rounds_roundReg_out[35]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_8_U3 ( .A0_t (Midori_rounds_roundReg_out[34]), .B0_t (Midori_rounds_roundReg_out[35]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_8_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n14), .Z0_t (Midori_rounds_SR_Result[19]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n13), .B0_t (Midori_rounds_roundReg_out[37]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n11), .Z0_t (Midori_rounds_SR_Result[17]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U16 ( .A0_t (Midori_rounds_roundReg_out[36]), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U15 ( .A0_t (Midori_rounds_roundReg_out[39]), .B0_t (Midori_rounds_roundReg_out[38]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U14 ( .A0_t (Midori_rounds_roundReg_out[38]), .B0_t (Midori_rounds_roundReg_out[39]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n7), .Z0_t (Midori_rounds_SR_Result[18]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n6), .B0_t (Midori_rounds_roundReg_out[37]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n5), .B0_t (Midori_rounds_roundReg_out[38]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U10 ( .A0_t (Midori_rounds_roundReg_out[36]), .B0_t (Midori_rounds_roundReg_out[39]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U9 ( .A0_t (Midori_rounds_roundReg_out[39]), .B0_t (Midori_rounds_roundReg_out[36]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_9_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n3), .Z0_t (Midori_rounds_SR_Result[16]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U7 ( .A0_t (Midori_rounds_roundReg_out[37]), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U6 ( .A0_t (Midori_rounds_roundReg_out[36]), .B0_t (Midori_rounds_sub_sBox_PRINCE_9_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U5 ( .A0_t (Midori_rounds_roundReg_out[38]), .B0_t (Midori_rounds_roundReg_out[39]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_9_U3 ( .A0_t (Midori_rounds_roundReg_out[38]), .B0_t (Midori_rounds_roundReg_out[39]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_9_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n14), .Z0_t (Midori_rounds_SR_Result[52]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U18 ( .A0_t (Midori_rounds_roundReg_out[41]), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U17 ( .A0_t (Midori_rounds_roundReg_out[40]), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U16 ( .A0_t (Midori_rounds_roundReg_out[42]), .B0_t (Midori_rounds_roundReg_out[43]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n9), .Z0_t (Midori_rounds_SR_Result[54]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n8), .B0_t (Midori_rounds_roundReg_out[41]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n7), .B0_t (Midori_rounds_roundReg_out[42]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U12 ( .A0_t (Midori_rounds_roundReg_out[40]), .B0_t (Midori_rounds_roundReg_out[43]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n5), .Z0_t (Midori_rounds_SR_Result[55]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U10 ( .A0_t (Midori_rounds_roundReg_out[41]), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U9 ( .A0_t (Midori_rounds_roundReg_out[42]), .B0_t (Midori_rounds_roundReg_out[43]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U8 ( .A0_t (Midori_rounds_roundReg_out[43]), .B0_t (Midori_rounds_roundReg_out[40]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_10_n2), .Z0_t (Midori_rounds_SR_Result[53]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_10_n1), .B0_t (Midori_rounds_roundReg_out[43]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U4 ( .A0_t (Midori_rounds_roundReg_out[42]), .B0_t (Midori_rounds_roundReg_out[40]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_10_U1 ( .A0_t (Midori_rounds_roundReg_out[42]), .B0_t (Midori_rounds_roundReg_out[40]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_10_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n14), .Z0_t (Midori_rounds_SR_Result[40]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U18 ( .A0_t (Midori_rounds_roundReg_out[45]), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U17 ( .A0_t (Midori_rounds_roundReg_out[44]), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U16 ( .A0_t (Midori_rounds_roundReg_out[46]), .B0_t (Midori_rounds_roundReg_out[47]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n9), .Z0_t (Midori_rounds_SR_Result[42]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n8), .B0_t (Midori_rounds_roundReg_out[45]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n7), .B0_t (Midori_rounds_roundReg_out[46]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U12 ( .A0_t (Midori_rounds_roundReg_out[44]), .B0_t (Midori_rounds_roundReg_out[47]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n5), .Z0_t (Midori_rounds_SR_Result[43]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U10 ( .A0_t (Midori_rounds_roundReg_out[45]), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U9 ( .A0_t (Midori_rounds_roundReg_out[46]), .B0_t (Midori_rounds_roundReg_out[47]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U8 ( .A0_t (Midori_rounds_roundReg_out[47]), .B0_t (Midori_rounds_roundReg_out[44]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_11_n2), .Z0_t (Midori_rounds_SR_Result[41]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_11_n1), .B0_t (Midori_rounds_roundReg_out[47]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U4 ( .A0_t (Midori_rounds_roundReg_out[46]), .B0_t (Midori_rounds_roundReg_out[44]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_11_U1 ( .A0_t (Midori_rounds_roundReg_out[46]), .B0_t (Midori_rounds_roundReg_out[44]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_11_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n14), .Z0_t (Midori_rounds_SR_Result[24]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U18 ( .A0_t (Midori_rounds_roundReg_out[49]), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U17 ( .A0_t (Midori_rounds_roundReg_out[48]), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U16 ( .A0_t (Midori_rounds_roundReg_out[50]), .B0_t (Midori_rounds_roundReg_out[51]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n9), .Z0_t (Midori_rounds_SR_Result[26]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n8), .B0_t (Midori_rounds_roundReg_out[49]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n7), .B0_t (Midori_rounds_roundReg_out[50]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U12 ( .A0_t (Midori_rounds_roundReg_out[48]), .B0_t (Midori_rounds_roundReg_out[51]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n5), .Z0_t (Midori_rounds_SR_Result[27]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U10 ( .A0_t (Midori_rounds_roundReg_out[49]), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U9 ( .A0_t (Midori_rounds_roundReg_out[50]), .B0_t (Midori_rounds_roundReg_out[51]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U8 ( .A0_t (Midori_rounds_roundReg_out[51]), .B0_t (Midori_rounds_roundReg_out[48]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_12_n2), .Z0_t (Midori_rounds_SR_Result[25]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_12_n1), .B0_t (Midori_rounds_roundReg_out[51]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U4 ( .A0_t (Midori_rounds_roundReg_out[50]), .B0_t (Midori_rounds_roundReg_out[48]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_12_U1 ( .A0_t (Midori_rounds_roundReg_out[50]), .B0_t (Midori_rounds_roundReg_out[48]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_12_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n14), .Z0_t (Midori_rounds_SR_Result[7]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n13), .B0_t (Midori_rounds_roundReg_out[53]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n11), .Z0_t (Midori_rounds_SR_Result[5]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U16 ( .A0_t (Midori_rounds_roundReg_out[52]), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U15 ( .A0_t (Midori_rounds_roundReg_out[55]), .B0_t (Midori_rounds_roundReg_out[54]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U14 ( .A0_t (Midori_rounds_roundReg_out[54]), .B0_t (Midori_rounds_roundReg_out[55]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n7), .Z0_t (Midori_rounds_SR_Result[6]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n6), .B0_t (Midori_rounds_roundReg_out[53]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n5), .B0_t (Midori_rounds_roundReg_out[54]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U10 ( .A0_t (Midori_rounds_roundReg_out[52]), .B0_t (Midori_rounds_roundReg_out[55]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U9 ( .A0_t (Midori_rounds_roundReg_out[55]), .B0_t (Midori_rounds_roundReg_out[52]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_13_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n3), .Z0_t (Midori_rounds_SR_Result[4]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U7 ( .A0_t (Midori_rounds_roundReg_out[53]), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U6 ( .A0_t (Midori_rounds_roundReg_out[52]), .B0_t (Midori_rounds_sub_sBox_PRINCE_13_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U5 ( .A0_t (Midori_rounds_roundReg_out[54]), .B0_t (Midori_rounds_roundReg_out[55]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_13_U3 ( .A0_t (Midori_rounds_roundReg_out[54]), .B0_t (Midori_rounds_roundReg_out[55]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_13_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n14), .Z0_t (Midori_rounds_SR_Result[35]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U18 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n13), .B0_t (Midori_rounds_roundReg_out[57]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U17 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n12), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n11), .Z0_t (Midori_rounds_SR_Result[33]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U16 ( .A0_t (Midori_rounds_roundReg_out[56]), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n10), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U15 ( .A0_t (Midori_rounds_roundReg_out[59]), .B0_t (Midori_rounds_roundReg_out[58]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U14 ( .A0_t (Midori_rounds_roundReg_out[58]), .B0_t (Midori_rounds_roundReg_out[59]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n12) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n7), .Z0_t (Midori_rounds_SR_Result[34]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U12 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n6), .B0_t (Midori_rounds_roundReg_out[57]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n5), .B0_t (Midori_rounds_roundReg_out[58]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n6) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U10 ( .A0_t (Midori_rounds_roundReg_out[56]), .B0_t (Midori_rounds_roundReg_out[59]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U9 ( .A0_t (Midori_rounds_roundReg_out[59]), .B0_t (Midori_rounds_roundReg_out[56]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U8 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_14_n13), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n3), .Z0_t (Midori_rounds_SR_Result[32]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U7 ( .A0_t (Midori_rounds_roundReg_out[57]), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n2), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n3) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U6 ( .A0_t (Midori_rounds_roundReg_out[56]), .B0_t (Midori_rounds_sub_sBox_PRINCE_14_n1), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U5 ( .A0_t (Midori_rounds_roundReg_out[58]), .B0_t (Midori_rounds_roundReg_out[59]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_14_U3 ( .A0_t (Midori_rounds_roundReg_out[58]), .B0_t (Midori_rounds_roundReg_out[59]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_14_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U19 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n15), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n14), .Z0_t (Midori_rounds_SR_Result[60]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U18 ( .A0_t (Midori_rounds_roundReg_out[61]), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n13), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n15) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U17 ( .A0_t (Midori_rounds_roundReg_out[60]), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n11), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n13) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U16 ( .A0_t (Midori_rounds_roundReg_out[62]), .B0_t (Midori_rounds_roundReg_out[63]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n11) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U15 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n10), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n9), .Z0_t (Midori_rounds_SR_Result[62]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U14 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n8), .B0_t (Midori_rounds_roundReg_out[61]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n10) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U13 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n7), .B0_t (Midori_rounds_roundReg_out[62]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n8) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U12 ( .A0_t (Midori_rounds_roundReg_out[60]), .B0_t (Midori_rounds_roundReg_out[63]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n7) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U11 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n9), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n5), .Z0_t (Midori_rounds_SR_Result[63]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U10 ( .A0_t (Midori_rounds_roundReg_out[61]), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n14), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n5) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U9 ( .A0_t (Midori_rounds_roundReg_out[62]), .B0_t (Midori_rounds_roundReg_out[63]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n14) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U8 ( .A0_t (Midori_rounds_roundReg_out[63]), .B0_t (Midori_rounds_roundReg_out[60]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n9) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U7 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n3), .B0_t (Midori_rounds_sub_sBox_PRINCE_15_n2), .Z0_t (Midori_rounds_SR_Result[61]) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U6 ( .A0_t (Midori_rounds_sub_sBox_PRINCE_15_n1), .B0_t (Midori_rounds_roundReg_out[63]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n2) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b1), .CB(1'b1), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U4 ( .A0_t (Midori_rounds_roundReg_out[62]), .B0_t (Midori_rounds_roundReg_out[60]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n1) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_sub_sBox_PRINCE_15_U1 ( .A0_t (Midori_rounds_roundReg_out[62]), .B0_t (Midori_rounds_roundReg_out[60]), .Z0_t (Midori_rounds_sub_sBox_PRINCE_15_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[0]), .B0_t (Midori_rounds_sub_ResultXORkey[0]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_0_U1_Y), .B0_t (Midori_rounds_SR_Result[0]), .Z0_t (Midori_rounds_mul_input[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[1]), .B0_t (Midori_rounds_sub_ResultXORkey[1]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_1_U1_Y), .B0_t (Midori_rounds_SR_Result[1]), .Z0_t (Midori_rounds_mul_input[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[2]), .B0_t (Midori_rounds_sub_ResultXORkey[2]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_2_U1_Y), .B0_t (Midori_rounds_SR_Result[2]), .Z0_t (Midori_rounds_mul_input[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[3]), .B0_t (Midori_rounds_sub_ResultXORkey[3]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_3_U1_Y), .B0_t (Midori_rounds_SR_Result[3]), .Z0_t (Midori_rounds_mul_input[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[4]), .B0_t (Midori_rounds_sub_ResultXORkey[4]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_4_U1_Y), .B0_t (Midori_rounds_SR_Result[4]), .Z0_t (Midori_rounds_mul_input[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[5]), .B0_t (Midori_rounds_sub_ResultXORkey[5]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_5_U1_Y), .B0_t (Midori_rounds_SR_Result[5]), .Z0_t (Midori_rounds_mul_input[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[6]), .B0_t (Midori_rounds_sub_ResultXORkey[6]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_6_U1_Y), .B0_t (Midori_rounds_SR_Result[6]), .Z0_t (Midori_rounds_mul_input[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[7]), .B0_t (Midori_rounds_sub_ResultXORkey[7]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_7_U1_Y), .B0_t (Midori_rounds_SR_Result[7]), .Z0_t (Midori_rounds_mul_input[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[8]), .B0_t (Midori_rounds_sub_ResultXORkey[8]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_8_U1_Y), .B0_t (Midori_rounds_SR_Result[8]), .Z0_t (Midori_rounds_mul_input[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[9]), .B0_t (Midori_rounds_sub_ResultXORkey[9]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_9_U1_Y), .B0_t (Midori_rounds_SR_Result[9]), .Z0_t (Midori_rounds_mul_input[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[10]), .B0_t (Midori_rounds_sub_ResultXORkey[10]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_10_U1_Y), .B0_t (Midori_rounds_SR_Result[10]), .Z0_t (Midori_rounds_mul_input[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[11]), .B0_t (Midori_rounds_sub_ResultXORkey[11]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_11_U1_Y), .B0_t (Midori_rounds_SR_Result[11]), .Z0_t (Midori_rounds_mul_input[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[12]), .B0_t (Midori_rounds_sub_ResultXORkey[12]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_12_U1_Y), .B0_t (Midori_rounds_SR_Result[12]), .Z0_t (Midori_rounds_mul_input[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[13]), .B0_t (Midori_rounds_sub_ResultXORkey[13]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_13_U1_Y), .B0_t (Midori_rounds_SR_Result[13]), .Z0_t (Midori_rounds_mul_input[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[14]), .B0_t (Midori_rounds_sub_ResultXORkey[14]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_14_U1_Y), .B0_t (Midori_rounds_SR_Result[14]), .Z0_t (Midori_rounds_mul_input[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[15]), .B0_t (Midori_rounds_sub_ResultXORkey[15]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_15_U1_Y), .B0_t (Midori_rounds_SR_Result[15]), .Z0_t (Midori_rounds_mul_input[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[16]), .B0_t (Midori_rounds_sub_ResultXORkey[16]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_16_U1_Y), .B0_t (Midori_rounds_SR_Result[16]), .Z0_t (Midori_rounds_mul_input[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[17]), .B0_t (Midori_rounds_sub_ResultXORkey[17]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_17_U1_Y), .B0_t (Midori_rounds_SR_Result[17]), .Z0_t (Midori_rounds_mul_input[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[18]), .B0_t (Midori_rounds_sub_ResultXORkey[18]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_18_U1_Y), .B0_t (Midori_rounds_SR_Result[18]), .Z0_t (Midori_rounds_mul_input[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[19]), .B0_t (Midori_rounds_sub_ResultXORkey[19]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_19_U1_Y), .B0_t (Midori_rounds_SR_Result[19]), .Z0_t (Midori_rounds_mul_input[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[20]), .B0_t (Midori_rounds_sub_ResultXORkey[20]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_20_U1_Y), .B0_t (Midori_rounds_SR_Result[20]), .Z0_t (Midori_rounds_mul_input[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[21]), .B0_t (Midori_rounds_sub_ResultXORkey[21]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_21_U1_Y), .B0_t (Midori_rounds_SR_Result[21]), .Z0_t (Midori_rounds_mul_input[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[22]), .B0_t (Midori_rounds_sub_ResultXORkey[22]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_22_U1_Y), .B0_t (Midori_rounds_SR_Result[22]), .Z0_t (Midori_rounds_mul_input[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[23]), .B0_t (Midori_rounds_sub_ResultXORkey[23]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_23_U1_Y), .B0_t (Midori_rounds_SR_Result[23]), .Z0_t (Midori_rounds_mul_input[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[24]), .B0_t (Midori_rounds_sub_ResultXORkey[24]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_24_U1_Y), .B0_t (Midori_rounds_SR_Result[24]), .Z0_t (Midori_rounds_mul_input[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[25]), .B0_t (Midori_rounds_sub_ResultXORkey[25]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_25_U1_Y), .B0_t (Midori_rounds_SR_Result[25]), .Z0_t (Midori_rounds_mul_input[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[26]), .B0_t (Midori_rounds_sub_ResultXORkey[26]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_26_U1_Y), .B0_t (Midori_rounds_SR_Result[26]), .Z0_t (Midori_rounds_mul_input[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[27]), .B0_t (Midori_rounds_sub_ResultXORkey[27]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_27_U1_Y), .B0_t (Midori_rounds_SR_Result[27]), .Z0_t (Midori_rounds_mul_input[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[28]), .B0_t (Midori_rounds_sub_ResultXORkey[28]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_28_U1_Y), .B0_t (Midori_rounds_SR_Result[28]), .Z0_t (Midori_rounds_mul_input[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[29]), .B0_t (Midori_rounds_sub_ResultXORkey[29]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_29_U1_Y), .B0_t (Midori_rounds_SR_Result[29]), .Z0_t (Midori_rounds_mul_input[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[30]), .B0_t (Midori_rounds_sub_ResultXORkey[30]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_30_U1_Y), .B0_t (Midori_rounds_SR_Result[30]), .Z0_t (Midori_rounds_mul_input[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[31]), .B0_t (Midori_rounds_sub_ResultXORkey[31]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_31_U1_Y), .B0_t (Midori_rounds_SR_Result[31]), .Z0_t (Midori_rounds_mul_input[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[32]), .B0_t (Midori_rounds_sub_ResultXORkey[32]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_32_U1_Y), .B0_t (Midori_rounds_SR_Result[32]), .Z0_t (Midori_rounds_mul_input[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[33]), .B0_t (Midori_rounds_sub_ResultXORkey[33]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_33_U1_Y), .B0_t (Midori_rounds_SR_Result[33]), .Z0_t (Midori_rounds_mul_input[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[34]), .B0_t (Midori_rounds_sub_ResultXORkey[34]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_34_U1_Y), .B0_t (Midori_rounds_SR_Result[34]), .Z0_t (Midori_rounds_mul_input[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[35]), .B0_t (Midori_rounds_sub_ResultXORkey[35]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_35_U1_Y), .B0_t (Midori_rounds_SR_Result[35]), .Z0_t (Midori_rounds_mul_input[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[36]), .B0_t (Midori_rounds_sub_ResultXORkey[36]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_36_U1_Y), .B0_t (Midori_rounds_SR_Result[36]), .Z0_t (Midori_rounds_mul_input[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[37]), .B0_t (Midori_rounds_sub_ResultXORkey[37]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_37_U1_Y), .B0_t (Midori_rounds_SR_Result[37]), .Z0_t (Midori_rounds_mul_input[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[38]), .B0_t (Midori_rounds_sub_ResultXORkey[38]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_38_U1_Y), .B0_t (Midori_rounds_SR_Result[38]), .Z0_t (Midori_rounds_mul_input[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[39]), .B0_t (Midori_rounds_sub_ResultXORkey[39]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_39_U1_Y), .B0_t (Midori_rounds_SR_Result[39]), .Z0_t (Midori_rounds_mul_input[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[40]), .B0_t (Midori_rounds_sub_ResultXORkey[40]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_40_U1_Y), .B0_t (Midori_rounds_SR_Result[40]), .Z0_t (Midori_rounds_mul_input[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[41]), .B0_t (Midori_rounds_sub_ResultXORkey[41]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_41_U1_Y), .B0_t (Midori_rounds_SR_Result[41]), .Z0_t (Midori_rounds_mul_input[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[42]), .B0_t (Midori_rounds_sub_ResultXORkey[42]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_42_U1_Y), .B0_t (Midori_rounds_SR_Result[42]), .Z0_t (Midori_rounds_mul_input[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[43]), .B0_t (Midori_rounds_sub_ResultXORkey[43]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_43_U1_Y), .B0_t (Midori_rounds_SR_Result[43]), .Z0_t (Midori_rounds_mul_input[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[44]), .B0_t (Midori_rounds_sub_ResultXORkey[44]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_44_U1_Y), .B0_t (Midori_rounds_SR_Result[44]), .Z0_t (Midori_rounds_mul_input[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[45]), .B0_t (Midori_rounds_sub_ResultXORkey[45]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_45_U1_Y), .B0_t (Midori_rounds_SR_Result[45]), .Z0_t (Midori_rounds_mul_input[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[46]), .B0_t (Midori_rounds_sub_ResultXORkey[46]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_46_U1_Y), .B0_t (Midori_rounds_SR_Result[46]), .Z0_t (Midori_rounds_mul_input[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[47]), .B0_t (Midori_rounds_sub_ResultXORkey[47]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_47_U1_Y), .B0_t (Midori_rounds_SR_Result[47]), .Z0_t (Midori_rounds_mul_input[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[48]), .B0_t (Midori_rounds_sub_ResultXORkey[48]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_48_U1_Y), .B0_t (Midori_rounds_SR_Result[48]), .Z0_t (Midori_rounds_mul_input[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[49]), .B0_t (Midori_rounds_sub_ResultXORkey[49]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_49_U1_Y), .B0_t (Midori_rounds_SR_Result[49]), .Z0_t (Midori_rounds_mul_input[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[50]), .B0_t (Midori_rounds_sub_ResultXORkey[50]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_50_U1_Y), .B0_t (Midori_rounds_SR_Result[50]), .Z0_t (Midori_rounds_mul_input[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[51]), .B0_t (Midori_rounds_sub_ResultXORkey[51]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_51_U1_Y), .B0_t (Midori_rounds_SR_Result[51]), .Z0_t (Midori_rounds_mul_input[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[52]), .B0_t (Midori_rounds_sub_ResultXORkey[52]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_52_U1_Y), .B0_t (Midori_rounds_SR_Result[52]), .Z0_t (Midori_rounds_mul_input[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[53]), .B0_t (Midori_rounds_sub_ResultXORkey[53]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_53_U1_Y), .B0_t (Midori_rounds_SR_Result[53]), .Z0_t (Midori_rounds_mul_input[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[54]), .B0_t (Midori_rounds_sub_ResultXORkey[54]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_54_U1_Y), .B0_t (Midori_rounds_SR_Result[54]), .Z0_t (Midori_rounds_mul_input[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[55]), .B0_t (Midori_rounds_sub_ResultXORkey[55]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_55_U1_Y), .B0_t (Midori_rounds_SR_Result[55]), .Z0_t (Midori_rounds_mul_input[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[56]), .B0_t (Midori_rounds_sub_ResultXORkey[56]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_56_U1_Y), .B0_t (Midori_rounds_SR_Result[56]), .Z0_t (Midori_rounds_mul_input[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[57]), .B0_t (Midori_rounds_sub_ResultXORkey[57]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_57_U1_Y), .B0_t (Midori_rounds_SR_Result[57]), .Z0_t (Midori_rounds_mul_input[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[58]), .B0_t (Midori_rounds_sub_ResultXORkey[58]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_58_U1_Y), .B0_t (Midori_rounds_SR_Result[58]), .Z0_t (Midori_rounds_mul_input[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[59]), .B0_t (Midori_rounds_sub_ResultXORkey[59]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_59_U1_Y), .B0_t (Midori_rounds_SR_Result[59]), .Z0_t (Midori_rounds_mul_input[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[60]), .B0_t (Midori_rounds_sub_ResultXORkey[60]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_60_U1_Y), .B0_t (Midori_rounds_SR_Result[60]), .Z0_t (Midori_rounds_mul_input[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[61]), .B0_t (Midori_rounds_sub_ResultXORkey[61]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_61_U1_Y), .B0_t (Midori_rounds_SR_Result[61]), .Z0_t (Midori_rounds_mul_input[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[62]), .B0_t (Midori_rounds_sub_ResultXORkey[62]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_62_U1_Y), .B0_t (Midori_rounds_SR_Result[62]), .Z0_t (Midori_rounds_mul_input[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_XOR1_U1 ( .A0_t (Midori_rounds_SR_Result[63]), .B0_t (Midori_rounds_sub_ResultXORkey[63]), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_X), .Z0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_mul_input_Inst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_mul_input_Inst_mux_inst_63_U1_Y), .B0_t (Midori_rounds_SR_Result[63]), .Z0_t (Midori_rounds_mul_input[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U24 ( .A0_t (Midori_rounds_mul_input[59]), .B0_t (Midori_rounds_mul_MC1_n8), .Z0_t (Midori_rounds_SR_Inv_Result[63]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U23 ( .A0_t (Midori_rounds_mul_input[63]), .B0_t (Midori_rounds_mul_MC1_n8), .Z0_t (Midori_rounds_SR_Inv_Result[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U22 ( .A0_t (Midori_rounds_mul_input[55]), .B0_t (Midori_rounds_mul_input[51]), .Z0_t (Midori_rounds_mul_MC1_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U21 ( .A0_t (Midori_rounds_mul_input[58]), .B0_t (Midori_rounds_mul_MC1_n7), .Z0_t (Midori_rounds_SR_Inv_Result[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U20 ( .A0_t (Midori_rounds_mul_input[62]), .B0_t (Midori_rounds_mul_MC1_n7), .Z0_t (Midori_rounds_SR_Inv_Result[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U19 ( .A0_t (Midori_rounds_mul_input[54]), .B0_t (Midori_rounds_mul_input[50]), .Z0_t (Midori_rounds_mul_MC1_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U18 ( .A0_t (Midori_rounds_mul_input[56]), .B0_t (Midori_rounds_mul_MC1_n6), .Z0_t (Midori_rounds_SR_Inv_Result[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U17 ( .A0_t (Midori_rounds_mul_input[60]), .B0_t (Midori_rounds_mul_MC1_n6), .Z0_t (Midori_rounds_SR_Inv_Result[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U16 ( .A0_t (Midori_rounds_mul_input[52]), .B0_t (Midori_rounds_mul_input[48]), .Z0_t (Midori_rounds_mul_MC1_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U15 ( .A0_t (Midori_rounds_mul_input[51]), .B0_t (Midori_rounds_mul_MC1_n5), .Z0_t (Midori_rounds_SR_Inv_Result[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U14 ( .A0_t (Midori_rounds_mul_input[55]), .B0_t (Midori_rounds_mul_MC1_n5), .Z0_t (Midori_rounds_SR_Inv_Result[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U13 ( .A0_t (Midori_rounds_mul_input[59]), .B0_t (Midori_rounds_mul_input[63]), .Z0_t (Midori_rounds_mul_MC1_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U12 ( .A0_t (Midori_rounds_mul_input[57]), .B0_t (Midori_rounds_mul_MC1_n4), .Z0_t (Midori_rounds_SR_Inv_Result[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U11 ( .A0_t (Midori_rounds_mul_input[61]), .B0_t (Midori_rounds_mul_MC1_n4), .Z0_t (Midori_rounds_SR_Inv_Result[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U10 ( .A0_t (Midori_rounds_mul_input[53]), .B0_t (Midori_rounds_mul_input[49]), .Z0_t (Midori_rounds_mul_MC1_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U9 ( .A0_t (Midori_rounds_mul_input[50]), .B0_t (Midori_rounds_mul_MC1_n3), .Z0_t (Midori_rounds_SR_Inv_Result[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U8 ( .A0_t (Midori_rounds_mul_input[54]), .B0_t (Midori_rounds_mul_MC1_n3), .Z0_t (Midori_rounds_SR_Inv_Result[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U7 ( .A0_t (Midori_rounds_mul_input[58]), .B0_t (Midori_rounds_mul_input[62]), .Z0_t (Midori_rounds_mul_MC1_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U6 ( .A0_t (Midori_rounds_mul_input[49]), .B0_t (Midori_rounds_mul_MC1_n2), .Z0_t (Midori_rounds_SR_Inv_Result[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U5 ( .A0_t (Midori_rounds_mul_input[53]), .B0_t (Midori_rounds_mul_MC1_n2), .Z0_t (Midori_rounds_SR_Inv_Result[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U4 ( .A0_t (Midori_rounds_mul_input[57]), .B0_t (Midori_rounds_mul_input[61]), .Z0_t (Midori_rounds_mul_MC1_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U3 ( .A0_t (Midori_rounds_mul_input[48]), .B0_t (Midori_rounds_mul_MC1_n1), .Z0_t (Midori_rounds_SR_Inv_Result[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U2 ( .A0_t (Midori_rounds_mul_input[52]), .B0_t (Midori_rounds_mul_MC1_n1), .Z0_t (Midori_rounds_SR_Inv_Result[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC1_U1 ( .A0_t (Midori_rounds_mul_input[56]), .B0_t (Midori_rounds_mul_input[60]), .Z0_t (Midori_rounds_mul_MC1_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U24 ( .A0_t (Midori_rounds_mul_input[43]), .B0_t (Midori_rounds_mul_MC2_n8), .Z0_t (Midori_rounds_SR_Inv_Result[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U23 ( .A0_t (Midori_rounds_mul_input[47]), .B0_t (Midori_rounds_mul_MC2_n8), .Z0_t (Midori_rounds_SR_Inv_Result[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U22 ( .A0_t (Midori_rounds_mul_input[39]), .B0_t (Midori_rounds_mul_input[35]), .Z0_t (Midori_rounds_mul_MC2_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U21 ( .A0_t (Midori_rounds_mul_input[42]), .B0_t (Midori_rounds_mul_MC2_n7), .Z0_t (Midori_rounds_SR_Inv_Result[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U20 ( .A0_t (Midori_rounds_mul_input[46]), .B0_t (Midori_rounds_mul_MC2_n7), .Z0_t (Midori_rounds_SR_Inv_Result[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U19 ( .A0_t (Midori_rounds_mul_input[38]), .B0_t (Midori_rounds_mul_input[34]), .Z0_t (Midori_rounds_mul_MC2_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U18 ( .A0_t (Midori_rounds_mul_input[40]), .B0_t (Midori_rounds_mul_MC2_n6), .Z0_t (Midori_rounds_SR_Inv_Result[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U17 ( .A0_t (Midori_rounds_mul_input[44]), .B0_t (Midori_rounds_mul_MC2_n6), .Z0_t (Midori_rounds_SR_Inv_Result[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U16 ( .A0_t (Midori_rounds_mul_input[36]), .B0_t (Midori_rounds_mul_input[32]), .Z0_t (Midori_rounds_mul_MC2_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U15 ( .A0_t (Midori_rounds_mul_input[35]), .B0_t (Midori_rounds_mul_MC2_n5), .Z0_t (Midori_rounds_SR_Inv_Result[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U14 ( .A0_t (Midori_rounds_mul_input[39]), .B0_t (Midori_rounds_mul_MC2_n5), .Z0_t (Midori_rounds_SR_Inv_Result[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U13 ( .A0_t (Midori_rounds_mul_input[43]), .B0_t (Midori_rounds_mul_input[47]), .Z0_t (Midori_rounds_mul_MC2_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U12 ( .A0_t (Midori_rounds_mul_input[41]), .B0_t (Midori_rounds_mul_MC2_n4), .Z0_t (Midori_rounds_SR_Inv_Result[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U11 ( .A0_t (Midori_rounds_mul_input[45]), .B0_t (Midori_rounds_mul_MC2_n4), .Z0_t (Midori_rounds_SR_Inv_Result[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U10 ( .A0_t (Midori_rounds_mul_input[37]), .B0_t (Midori_rounds_mul_input[33]), .Z0_t (Midori_rounds_mul_MC2_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U9 ( .A0_t (Midori_rounds_mul_input[34]), .B0_t (Midori_rounds_mul_MC2_n3), .Z0_t (Midori_rounds_SR_Inv_Result[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U8 ( .A0_t (Midori_rounds_mul_input[38]), .B0_t (Midori_rounds_mul_MC2_n3), .Z0_t (Midori_rounds_SR_Inv_Result[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U7 ( .A0_t (Midori_rounds_mul_input[42]), .B0_t (Midori_rounds_mul_input[46]), .Z0_t (Midori_rounds_mul_MC2_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U6 ( .A0_t (Midori_rounds_mul_input[33]), .B0_t (Midori_rounds_mul_MC2_n2), .Z0_t (Midori_rounds_SR_Inv_Result[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U5 ( .A0_t (Midori_rounds_mul_input[37]), .B0_t (Midori_rounds_mul_MC2_n2), .Z0_t (Midori_rounds_SR_Inv_Result[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U4 ( .A0_t (Midori_rounds_mul_input[41]), .B0_t (Midori_rounds_mul_input[45]), .Z0_t (Midori_rounds_mul_MC2_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U3 ( .A0_t (Midori_rounds_mul_input[32]), .B0_t (Midori_rounds_mul_MC2_n1), .Z0_t (Midori_rounds_SR_Inv_Result[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U2 ( .A0_t (Midori_rounds_mul_input[36]), .B0_t (Midori_rounds_mul_MC2_n1), .Z0_t (Midori_rounds_SR_Inv_Result[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC2_U1 ( .A0_t (Midori_rounds_mul_input[40]), .B0_t (Midori_rounds_mul_input[44]), .Z0_t (Midori_rounds_mul_MC2_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U24 ( .A0_t (Midori_rounds_mul_input[27]), .B0_t (Midori_rounds_mul_MC3_n8), .Z0_t (Midori_rounds_SR_Inv_Result[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U23 ( .A0_t (Midori_rounds_mul_input[31]), .B0_t (Midori_rounds_mul_MC3_n8), .Z0_t (Midori_rounds_SR_Inv_Result[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U22 ( .A0_t (Midori_rounds_mul_input[23]), .B0_t (Midori_rounds_mul_input[19]), .Z0_t (Midori_rounds_mul_MC3_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U21 ( .A0_t (Midori_rounds_mul_input[26]), .B0_t (Midori_rounds_mul_MC3_n7), .Z0_t (Midori_rounds_SR_Inv_Result[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U20 ( .A0_t (Midori_rounds_mul_input[30]), .B0_t (Midori_rounds_mul_MC3_n7), .Z0_t (Midori_rounds_SR_Inv_Result[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U19 ( .A0_t (Midori_rounds_mul_input[22]), .B0_t (Midori_rounds_mul_input[18]), .Z0_t (Midori_rounds_mul_MC3_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U18 ( .A0_t (Midori_rounds_mul_input[24]), .B0_t (Midori_rounds_mul_MC3_n6), .Z0_t (Midori_rounds_SR_Inv_Result[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U17 ( .A0_t (Midori_rounds_mul_input[28]), .B0_t (Midori_rounds_mul_MC3_n6), .Z0_t (Midori_rounds_SR_Inv_Result[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U16 ( .A0_t (Midori_rounds_mul_input[20]), .B0_t (Midori_rounds_mul_input[16]), .Z0_t (Midori_rounds_mul_MC3_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U15 ( .A0_t (Midori_rounds_mul_input[19]), .B0_t (Midori_rounds_mul_MC3_n5), .Z0_t (Midori_rounds_SR_Inv_Result[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U14 ( .A0_t (Midori_rounds_mul_input[23]), .B0_t (Midori_rounds_mul_MC3_n5), .Z0_t (Midori_rounds_SR_Inv_Result[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U13 ( .A0_t (Midori_rounds_mul_input[27]), .B0_t (Midori_rounds_mul_input[31]), .Z0_t (Midori_rounds_mul_MC3_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U12 ( .A0_t (Midori_rounds_mul_input[25]), .B0_t (Midori_rounds_mul_MC3_n4), .Z0_t (Midori_rounds_SR_Inv_Result[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U11 ( .A0_t (Midori_rounds_mul_input[29]), .B0_t (Midori_rounds_mul_MC3_n4), .Z0_t (Midori_rounds_SR_Inv_Result[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U10 ( .A0_t (Midori_rounds_mul_input[21]), .B0_t (Midori_rounds_mul_input[17]), .Z0_t (Midori_rounds_mul_MC3_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U9 ( .A0_t (Midori_rounds_mul_input[18]), .B0_t (Midori_rounds_mul_MC3_n3), .Z0_t (Midori_rounds_SR_Inv_Result[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U8 ( .A0_t (Midori_rounds_mul_input[22]), .B0_t (Midori_rounds_mul_MC3_n3), .Z0_t (Midori_rounds_SR_Inv_Result[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U7 ( .A0_t (Midori_rounds_mul_input[26]), .B0_t (Midori_rounds_mul_input[30]), .Z0_t (Midori_rounds_mul_MC3_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U6 ( .A0_t (Midori_rounds_mul_input[17]), .B0_t (Midori_rounds_mul_MC3_n2), .Z0_t (Midori_rounds_SR_Inv_Result[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U5 ( .A0_t (Midori_rounds_mul_input[21]), .B0_t (Midori_rounds_mul_MC3_n2), .Z0_t (Midori_rounds_SR_Inv_Result[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U4 ( .A0_t (Midori_rounds_mul_input[25]), .B0_t (Midori_rounds_mul_input[29]), .Z0_t (Midori_rounds_mul_MC3_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U3 ( .A0_t (Midori_rounds_mul_input[16]), .B0_t (Midori_rounds_mul_MC3_n1), .Z0_t (Midori_rounds_SR_Inv_Result[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U2 ( .A0_t (Midori_rounds_mul_input[20]), .B0_t (Midori_rounds_mul_MC3_n1), .Z0_t (Midori_rounds_SR_Inv_Result[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC3_U1 ( .A0_t (Midori_rounds_mul_input[24]), .B0_t (Midori_rounds_mul_input[28]), .Z0_t (Midori_rounds_mul_MC3_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U24 ( .A0_t (Midori_rounds_mul_input[11]), .B0_t (Midori_rounds_mul_MC4_n8), .Z0_t (Midori_rounds_SR_Inv_Result[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U23 ( .A0_t (Midori_rounds_mul_input[15]), .B0_t (Midori_rounds_mul_MC4_n8), .Z0_t (Midori_rounds_SR_Inv_Result[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U22 ( .A0_t (Midori_rounds_mul_input[7]), .B0_t (Midori_rounds_mul_input[3]), .Z0_t (Midori_rounds_mul_MC4_n8) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U21 ( .A0_t (Midori_rounds_mul_input[10]), .B0_t (Midori_rounds_mul_MC4_n7), .Z0_t (Midori_rounds_SR_Inv_Result[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U20 ( .A0_t (Midori_rounds_mul_input[14]), .B0_t (Midori_rounds_mul_MC4_n7), .Z0_t (Midori_rounds_SR_Inv_Result[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U19 ( .A0_t (Midori_rounds_mul_input[6]), .B0_t (Midori_rounds_mul_input[2]), .Z0_t (Midori_rounds_mul_MC4_n7) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U18 ( .A0_t (Midori_rounds_mul_input[8]), .B0_t (Midori_rounds_mul_MC4_n6), .Z0_t (Midori_rounds_SR_Inv_Result[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U17 ( .A0_t (Midori_rounds_mul_input[12]), .B0_t (Midori_rounds_mul_MC4_n6), .Z0_t (Midori_rounds_SR_Inv_Result[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U16 ( .A0_t (Midori_rounds_mul_input[4]), .B0_t (Midori_rounds_mul_input[0]), .Z0_t (Midori_rounds_mul_MC4_n6) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U15 ( .A0_t (Midori_rounds_mul_input[3]), .B0_t (Midori_rounds_mul_MC4_n5), .Z0_t (Midori_rounds_SR_Inv_Result[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U14 ( .A0_t (Midori_rounds_mul_input[7]), .B0_t (Midori_rounds_mul_MC4_n5), .Z0_t (Midori_rounds_SR_Inv_Result[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U13 ( .A0_t (Midori_rounds_mul_input[11]), .B0_t (Midori_rounds_mul_input[15]), .Z0_t (Midori_rounds_mul_MC4_n5) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U12 ( .A0_t (Midori_rounds_mul_input[9]), .B0_t (Midori_rounds_mul_MC4_n4), .Z0_t (Midori_rounds_SR_Inv_Result[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U11 ( .A0_t (Midori_rounds_mul_input[13]), .B0_t (Midori_rounds_mul_MC4_n4), .Z0_t (Midori_rounds_SR_Inv_Result[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U10 ( .A0_t (Midori_rounds_mul_input[5]), .B0_t (Midori_rounds_mul_input[1]), .Z0_t (Midori_rounds_mul_MC4_n4) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U9 ( .A0_t (Midori_rounds_mul_input[2]), .B0_t (Midori_rounds_mul_MC4_n3), .Z0_t (Midori_rounds_SR_Inv_Result[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U8 ( .A0_t (Midori_rounds_mul_input[6]), .B0_t (Midori_rounds_mul_MC4_n3), .Z0_t (Midori_rounds_SR_Inv_Result[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U7 ( .A0_t (Midori_rounds_mul_input[10]), .B0_t (Midori_rounds_mul_input[14]), .Z0_t (Midori_rounds_mul_MC4_n3) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U6 ( .A0_t (Midori_rounds_mul_input[1]), .B0_t (Midori_rounds_mul_MC4_n2), .Z0_t (Midori_rounds_SR_Inv_Result[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U5 ( .A0_t (Midori_rounds_mul_input[5]), .B0_t (Midori_rounds_mul_MC4_n2), .Z0_t (Midori_rounds_SR_Inv_Result[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U4 ( .A0_t (Midori_rounds_mul_input[9]), .B0_t (Midori_rounds_mul_input[13]), .Z0_t (Midori_rounds_mul_MC4_n2) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U3 ( .A0_t (Midori_rounds_mul_input[0]), .B0_t (Midori_rounds_mul_MC4_n1), .Z0_t (Midori_rounds_SR_Inv_Result[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U2 ( .A0_t (Midori_rounds_mul_input[4]), .B0_t (Midori_rounds_mul_MC4_n1), .Z0_t (Midori_rounds_SR_Inv_Result[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b1), .FF(1'b0)) Midori_rounds_mul_MC4_U1 ( .A0_t (Midori_rounds_mul_input[8]), .B0_t (Midori_rounds_mul_input[12]), .Z0_t (Midori_rounds_mul_MC4_n1) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[0]), .B0_t (Midori_rounds_SR_Inv_Result[0]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_0_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_0_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[0]), .Z0_t (Midori_rounds_round_Result[0]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[1]), .B0_t (Midori_rounds_SR_Inv_Result[1]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_1_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_1_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[1]), .Z0_t (Midori_rounds_round_Result[1]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[2]), .B0_t (Midori_rounds_SR_Inv_Result[2]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_2_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_2_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[2]), .Z0_t (Midori_rounds_round_Result[2]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[3]), .B0_t (Midori_rounds_SR_Inv_Result[3]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_3_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_3_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[3]), .Z0_t (Midori_rounds_round_Result[3]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[4]), .B0_t (Midori_rounds_SR_Inv_Result[4]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_4_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_4_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[4]), .Z0_t (Midori_rounds_round_Result[4]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[5]), .B0_t (Midori_rounds_SR_Inv_Result[5]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_5_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_5_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[5]), .Z0_t (Midori_rounds_round_Result[5]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[6]), .B0_t (Midori_rounds_SR_Inv_Result[6]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_6_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_6_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[6]), .Z0_t (Midori_rounds_round_Result[6]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[7]), .B0_t (Midori_rounds_SR_Inv_Result[7]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_7_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_7_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[7]), .Z0_t (Midori_rounds_round_Result[7]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[8]), .B0_t (Midori_rounds_SR_Inv_Result[8]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_8_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_8_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[8]), .Z0_t (Midori_rounds_round_Result[8]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[9]), .B0_t (Midori_rounds_SR_Inv_Result[9]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_9_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_9_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[9]), .Z0_t (Midori_rounds_round_Result[9]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[10]), .B0_t (Midori_rounds_SR_Inv_Result[10]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_10_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_10_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[10]), .Z0_t (Midori_rounds_round_Result[10]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[11]), .B0_t (Midori_rounds_SR_Inv_Result[11]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_11_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_11_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[11]), .Z0_t (Midori_rounds_round_Result[11]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[12]), .B0_t (Midori_rounds_SR_Inv_Result[12]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_12_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_12_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[12]), .Z0_t (Midori_rounds_round_Result[12]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[13]), .B0_t (Midori_rounds_SR_Inv_Result[13]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_13_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_13_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[13]), .Z0_t (Midori_rounds_round_Result[13]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[14]), .B0_t (Midori_rounds_SR_Inv_Result[14]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_14_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_14_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[14]), .Z0_t (Midori_rounds_round_Result[14]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[15]), .B0_t (Midori_rounds_SR_Inv_Result[15]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_15_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_15_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[15]), .Z0_t (Midori_rounds_round_Result[15]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[16]), .B0_t (Midori_rounds_SR_Inv_Result[16]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_16_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_16_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[16]), .Z0_t (Midori_rounds_round_Result[16]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[17]), .B0_t (Midori_rounds_SR_Inv_Result[17]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_17_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_17_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[17]), .Z0_t (Midori_rounds_round_Result[17]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[18]), .B0_t (Midori_rounds_SR_Inv_Result[18]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_18_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_18_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[18]), .Z0_t (Midori_rounds_round_Result[18]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[19]), .B0_t (Midori_rounds_SR_Inv_Result[19]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_19_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_19_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[19]), .Z0_t (Midori_rounds_round_Result[19]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[20]), .B0_t (Midori_rounds_SR_Inv_Result[20]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_20_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_20_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[20]), .Z0_t (Midori_rounds_round_Result[20]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[21]), .B0_t (Midori_rounds_SR_Inv_Result[21]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_21_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_21_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[21]), .Z0_t (Midori_rounds_round_Result[21]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[22]), .B0_t (Midori_rounds_SR_Inv_Result[22]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_22_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_22_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[22]), .Z0_t (Midori_rounds_round_Result[22]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[23]), .B0_t (Midori_rounds_SR_Inv_Result[23]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_23_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_23_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[23]), .Z0_t (Midori_rounds_round_Result[23]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[24]), .B0_t (Midori_rounds_SR_Inv_Result[24]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_24_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_24_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[24]), .Z0_t (Midori_rounds_round_Result[24]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[25]), .B0_t (Midori_rounds_SR_Inv_Result[25]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_25_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_25_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[25]), .Z0_t (Midori_rounds_round_Result[25]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[26]), .B0_t (Midori_rounds_SR_Inv_Result[26]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_26_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_26_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[26]), .Z0_t (Midori_rounds_round_Result[26]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[27]), .B0_t (Midori_rounds_SR_Inv_Result[27]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_27_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_27_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[27]), .Z0_t (Midori_rounds_round_Result[27]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[28]), .B0_t (Midori_rounds_SR_Inv_Result[28]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_28_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_28_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[28]), .Z0_t (Midori_rounds_round_Result[28]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[29]), .B0_t (Midori_rounds_SR_Inv_Result[29]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_29_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_29_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[29]), .Z0_t (Midori_rounds_round_Result[29]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[30]), .B0_t (Midori_rounds_SR_Inv_Result[30]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_30_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_30_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[30]), .Z0_t (Midori_rounds_round_Result[30]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[31]), .B0_t (Midori_rounds_SR_Inv_Result[31]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_31_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_31_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[31]), .Z0_t (Midori_rounds_round_Result[31]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[32]), .B0_t (Midori_rounds_SR_Inv_Result[32]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_32_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_32_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[32]), .Z0_t (Midori_rounds_round_Result[32]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[33]), .B0_t (Midori_rounds_SR_Inv_Result[33]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_33_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_33_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[33]), .Z0_t (Midori_rounds_round_Result[33]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[34]), .B0_t (Midori_rounds_SR_Inv_Result[34]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_34_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_34_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[34]), .Z0_t (Midori_rounds_round_Result[34]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[35]), .B0_t (Midori_rounds_SR_Inv_Result[35]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_35_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_35_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[35]), .Z0_t (Midori_rounds_round_Result[35]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[36]), .B0_t (Midori_rounds_SR_Inv_Result[36]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_36_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_36_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[36]), .Z0_t (Midori_rounds_round_Result[36]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[37]), .B0_t (Midori_rounds_SR_Inv_Result[37]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_37_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_37_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[37]), .Z0_t (Midori_rounds_round_Result[37]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[38]), .B0_t (Midori_rounds_SR_Inv_Result[38]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_38_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_38_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[38]), .Z0_t (Midori_rounds_round_Result[38]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[39]), .B0_t (Midori_rounds_SR_Inv_Result[39]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_39_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_39_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[39]), .Z0_t (Midori_rounds_round_Result[39]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[40]), .B0_t (Midori_rounds_SR_Inv_Result[40]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_40_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_40_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[40]), .Z0_t (Midori_rounds_round_Result[40]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[41]), .B0_t (Midori_rounds_SR_Inv_Result[41]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_41_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_41_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[41]), .Z0_t (Midori_rounds_round_Result[41]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[42]), .B0_t (Midori_rounds_SR_Inv_Result[42]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_42_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_42_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[42]), .Z0_t (Midori_rounds_round_Result[42]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[43]), .B0_t (Midori_rounds_SR_Inv_Result[43]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_43_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_43_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[43]), .Z0_t (Midori_rounds_round_Result[43]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[44]), .B0_t (Midori_rounds_SR_Inv_Result[44]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_44_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_44_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[44]), .Z0_t (Midori_rounds_round_Result[44]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[45]), .B0_t (Midori_rounds_SR_Inv_Result[45]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_45_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_45_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[45]), .Z0_t (Midori_rounds_round_Result[45]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[46]), .B0_t (Midori_rounds_SR_Inv_Result[46]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_46_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_46_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[46]), .Z0_t (Midori_rounds_round_Result[46]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[47]), .B0_t (Midori_rounds_SR_Inv_Result[47]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_47_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_47_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[47]), .Z0_t (Midori_rounds_round_Result[47]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[48]), .B0_t (Midori_rounds_SR_Inv_Result[48]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_48_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_48_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[48]), .Z0_t (Midori_rounds_round_Result[48]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[49]), .B0_t (Midori_rounds_SR_Inv_Result[49]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_49_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_49_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[49]), .Z0_t (Midori_rounds_round_Result[49]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[50]), .B0_t (Midori_rounds_SR_Inv_Result[50]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_50_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_50_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[50]), .Z0_t (Midori_rounds_round_Result[50]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[51]), .B0_t (Midori_rounds_SR_Inv_Result[51]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_51_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_51_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[51]), .Z0_t (Midori_rounds_round_Result[51]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[52]), .B0_t (Midori_rounds_SR_Inv_Result[52]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_52_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_52_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[52]), .Z0_t (Midori_rounds_round_Result[52]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[53]), .B0_t (Midori_rounds_SR_Inv_Result[53]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_53_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_53_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[53]), .Z0_t (Midori_rounds_round_Result[53]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[54]), .B0_t (Midori_rounds_SR_Inv_Result[54]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_54_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_54_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[54]), .Z0_t (Midori_rounds_round_Result[54]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[55]), .B0_t (Midori_rounds_SR_Inv_Result[55]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_55_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_55_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[55]), .Z0_t (Midori_rounds_round_Result[55]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[56]), .B0_t (Midori_rounds_SR_Inv_Result[56]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_56_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_56_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[56]), .Z0_t (Midori_rounds_round_Result[56]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[57]), .B0_t (Midori_rounds_SR_Inv_Result[57]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_57_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_57_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[57]), .Z0_t (Midori_rounds_round_Result[57]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[58]), .B0_t (Midori_rounds_SR_Inv_Result[58]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_58_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_58_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[58]), .Z0_t (Midori_rounds_round_Result[58]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[59]), .B0_t (Midori_rounds_SR_Inv_Result[59]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_59_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_59_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[59]), .Z0_t (Midori_rounds_round_Result[59]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[60]), .B0_t (Midori_rounds_SR_Inv_Result[60]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_60_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_60_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[60]), .Z0_t (Midori_rounds_round_Result[60]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[61]), .B0_t (Midori_rounds_SR_Inv_Result[61]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_61_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_61_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[61]), .Z0_t (Midori_rounds_round_Result[61]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[62]), .B0_t (Midori_rounds_SR_Inv_Result[62]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_62_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_62_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[62]), .Z0_t (Midori_rounds_round_Result[62]) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_XOR1_U1 ( .A0_t (Midori_rounds_mul_ResultXORkey[63]), .B0_t (Midori_rounds_SR_Inv_Result[63]), .Z0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_X) ) ;
    (* Keep *) nonlinear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_AND1_U1 ( .A0_t (enc_dec), .B0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_X), .Z0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_Y) ) ;
    (* Keep *) linear_LMDPL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b0)) Midori_rounds_Res_Inst_mux_inst_63_U1_XOR2_U1 ( .A0_t (Midori_rounds_Res_Inst_mux_inst_63_U1_Y), .B0_t (Midori_rounds_mul_ResultXORkey[63]), .Z0_t (Midori_rounds_round_Result[63]) ) ;
    (* Keep *) combined_WDDL_primitive #(.CA(1'b0), .CB(1'b0), .CZ(1'b0), .FF(1'b1), .NL(1'b0)) new_AGEMA_gate_1804 ( .A0_t (controller_roundCounter_N7), .B0_t (1'b0), .Z0_t (round_Signal[0]) ) ;

    /* register cells */
endmodule
